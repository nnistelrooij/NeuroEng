module run_network
#(
	parameter WIDTH = 8,
	parameter HEIGHT = 7,
	parameter NUM_POS_WEIGHTS = 3,
	parameter bit [WIDTH:0] WEIGHTS [0:HEIGHT - 1] = '{9'd60, 9'd60, 9'd60, 9'd60, 9'd60, 9'd60, 9'd60}
)
(
	input wire clk,  // clock signal
	input wire [HEIGHT - 1:0] pixels,  // binary inputs
	input wire start,  // active high start signal
	// binary outputs; 00: don't know, 01: pos class, 10: neg class
	output wire [1:0] neuron_out,
	output [$clog2(HEIGHT * (2 ** WIDTH - 1) + 1) - 1:0] balance_out
);
	reg running = 0;  // whether network is running
	// number of iterations network has been running
	reg [$clog2(HEIGHT * (2 **(WIDTH + 1) + 2)) - 1:0] iters = 0;

	network #(.WIDTH(WIDTH), .HEIGHT(HEIGHT), .NUM_POS_WEIGHTS(NUM_POS_WEIGHTS), .WEIGHTS(WEIGHTS)) N (
		.clk(running & clk),
		.rst(!start),
		.pixels(pixels),
		.neuron_out(neuron_out[0]),
		.balance_out(balance_out)
	);
	
	always @(posedge clk, posedge start) begin
		if (start) begin
			running = 1;
			iters = 0;
		end else if (iters == (HEIGHT * (2 **(WIDTH + 1) + 2) - 1)) begin
			running = 0;
			iters = 0;
		end else begin
			iters = iters + running;
		end
	end
	
	assign neuron_out[1] = !start & !running & !neuron_out[0];
endmodule

module test_all_images;
	reg clk = 0;
	reg [783:0] pixels = 0;
	reg start = 0;
	wire [1:0] neuron_out;
	reg [1:0] expected_neuron_out = 0;
	reg [$clog2(1038) - 1:0] guessed_neuron_out = 0;

	run_network #(
		.WIDTH(8),
		.HEIGHT(784),
		.WEIGHTS('{9'd0,9'd260,9'd261,9'd7,9'd0,9'd258,9'd0,9'd273,9'd261,9'd266,9'd2,9'd258,9'd6,9'd2,9'd264,9'd1,9'd260,9'd0,9'd1,9'd260,9'd5,9'd1,9'd0,9'd265,9'd259,9'd260,9'd6,9'd15,9'd0,9'd270,9'd264,9'd5,9'd262,9'd17,9'd266,9'd5,9'd0,9'd259,9'd258,9'd259,9'd4,9'd261,9'd0,9'd261,9'd11,9'd6,9'd1,9'd258,9'd260,9'd3,9'd258,9'd0,9'd260,9'd6,9'd3,9'd1,9'd5,9'd258,9'd258,9'd5,9'd0,9'd3,9'd0,9'd0,9'd266,9'd0,9'd265,9'd264,9'd261,9'd12,9'd4,9'd0,9'd292,9'd288,9'd259,9'd264,9'd0,9'd5,9'd0,9'd3,9'd7,9'd5,9'd258,9'd2,9'd1,9'd1,9'd3,9'd5,9'd264,9'd0,9'd261,9'd257,9'd294,9'd259,9'd305,9'd310,9'd347,9'd281,9'd293,9'd349,9'd330,9'd312,9'd322,9'd267,9'd268,9'd262,9'd4,9'd259,9'd4,9'd261,9'd264,9'd11,9'd257,9'd18,9'd6,9'd2,9'd2,9'd273,9'd268,9'd323,9'd297,9'd332,9'd389,9'd471,9'd509,9'd507,9'd419,9'd473,9'd475,9'd382,9'd399,9'd351,9'd286,9'd277,9'd6,9'd261,9'd8,9'd270,9'd1,9'd7,9'd0,9'd261,9'd0,9'd264,9'd261,9'd40,9'd32,9'd306,9'd35,9'd109,9'd274,9'd291,9'd305,9'd305,9'd10,9'd280,9'd285,9'd345,9'd389,9'd393,9'd436,9'd401,9'd358,9'd344,9'd8,9'd266,9'd257,9'd0,9'd258,9'd259,9'd272,9'd8,9'd75,9'd152,9'd78,9'd262,9'd92,9'd337,9'd268,9'd335,9'd38,9'd43,9'd19,9'd327,9'd305,9'd81,9'd336,9'd327,9'd341,9'd267,9'd56,9'd319,9'd275,9'd0,9'd5,9'd0,9'd266,9'd0,9'd0,9'd58,9'd149,9'd264,9'd17,9'd124,9'd359,9'd120,9'd37,9'd48,9'd310,9'd259,9'd298,9'd26,9'd286,9'd39,9'd85,9'd265,9'd119,9'd39,9'd82,9'd68,9'd331,9'd0,9'd7,9'd12,9'd260,9'd17,9'd52,9'd22,9'd78,9'd0,9'd111,9'd78,9'd62,9'd91,9'd303,9'd271,9'd102,9'd317,9'd29,9'd261,9'd275,9'd86,9'd276,9'd53,9'd271,9'd78,9'd18,9'd68,9'd287,9'd1,9'd4,9'd3,9'd3,9'd10,9'd35,9'd88,9'd107,9'd279,9'd51,9'd26,9'd13,9'd0,9'd327,9'd260,9'd46,9'd53,9'd296,9'd12,9'd31,9'd278,9'd34,9'd60,9'd358,9'd58,9'd23,9'd2,9'd17,9'd3,9'd22,9'd26,9'd8,9'd23,9'd40,9'd15,9'd95,9'd48,9'd68,9'd18,9'd1,9'd136,9'd0,9'd45,9'd285,9'd305,9'd46,9'd120,9'd105,9'd261,9'd55,9'd91,9'd305,9'd37,9'd112,9'd269,9'd25,9'd24,9'd26,9'd6,9'd258,9'd27,9'd76,9'd112,9'd78,9'd261,9'd101,9'd39,9'd57,9'd264,9'd187,9'd95,9'd0,9'd273,9'd104,9'd61,9'd149,9'd141,9'd85,9'd291,9'd78,9'd66,9'd114,9'd57,9'd58,9'd6,9'd267,9'd8,9'd257,9'd17,9'd73,9'd79,9'd56,9'd131,9'd77,9'd117,9'd233,9'd267,9'd328,9'd323,9'd426,9'd280,9'd304,9'd2,9'd30,9'd263,9'd56,9'd308,9'd336,9'd104,9'd109,9'd292,9'd76,9'd0,9'd11,9'd259,9'd259,9'd9,9'd30,9'd54,9'd48,9'd101,9'd299,9'd263,9'd298,9'd98,9'd118,9'd316,9'd504,9'd436,9'd337,9'd95,9'd286,9'd309,9'd282,9'd281,9'd56,9'd92,9'd101,9'd55,9'd25,9'd268,9'd4,9'd10,9'd4,9'd3,9'd11,9'd25,9'd42,9'd72,9'd28,9'd116,9'd20,9'd96,9'd73,9'd276,9'd355,9'd314,9'd296,9'd363,9'd302,9'd83,9'd64,9'd96,9'd54,9'd348,9'd86,9'd9,9'd20,9'd0,9'd0,9'd267,9'd266,9'd2,9'd257,9'd69,9'd11,9'd263,9'd47,9'd55,9'd19,9'd307,9'd101,9'd60,9'd374,9'd318,9'd330,9'd34,9'd288,9'd32,9'd57,9'd26,9'd301,9'd23,9'd56,9'd294,9'd313,9'd7,9'd261,9'd4,9'd0,9'd258,9'd266,9'd270,9'd5,9'd50,9'd133,9'd68,9'd70,9'd264,9'd278,9'd273,9'd340,9'd363,9'd51,9'd46,9'd135,9'd70,9'd271,9'd274,9'd333,9'd264,9'd324,9'd351,9'd324,9'd0,9'd0,9'd0,9'd6,9'd257,9'd263,9'd354,9'd343,9'd377,9'd21,9'd0,9'd296,9'd45,9'd312,9'd33,9'd298,9'd96,9'd121,9'd100,9'd147,9'd348,9'd267,9'd331,9'd265,9'd0,9'd273,9'd278,9'd79,9'd25,9'd257,9'd262,9'd6,9'd5,9'd263,9'd351,9'd391,9'd365,9'd401,9'd384,9'd296,9'd294,9'd329,9'd1,9'd306,9'd45,9'd53,9'd306,9'd395,9'd330,9'd96,9'd372,9'd57,9'd291,9'd312,9'd85,9'd73,9'd1,9'd265,9'd1,9'd7,9'd264,9'd261,9'd321,9'd370,9'd476,9'd352,9'd4,9'd26,9'd308,9'd78,9'd255,9'd302,9'd306,9'd282,9'd328,9'd283,9'd265,9'd333,9'd332,9'd294,9'd327,9'd357,9'd87,9'd120,9'd259,9'd261,9'd262,9'd259,9'd1,9'd265,9'd319,9'd449,9'd407,9'd381,9'd352,9'd284,9'd322,9'd53,9'd112,9'd88,9'd16,9'd306,9'd312,9'd283,9'd362,9'd404,9'd372,9'd397,9'd428,9'd472,9'd10,9'd52,9'd263,9'd261,9'd263,9'd257,9'd7,9'd319,9'd367,9'd407,9'd410,9'd321,9'd456,9'd351,9'd35,9'd260,9'd123,9'd108,9'd8,9'd326,9'd325,9'd364,9'd310,9'd449,9'd378,9'd415,9'd340,9'd409,9'd304,9'd259,9'd3,9'd260,9'd0,9'd0,9'd258,9'd277,9'd369,9'd395,9'd106,9'd289,9'd345,9'd351,9'd302,9'd446,9'd385,9'd42,9'd27,9'd285,9'd31,9'd359,9'd379,9'd343,9'd299,9'd365,9'd363,9'd365,9'd289,9'd11,9'd0,9'd4,9'd1,9'd9,9'd257,9'd4,9'd342,9'd295,9'd308,9'd31,9'd36,9'd389,9'd285,9'd302,9'd364,9'd257,9'd263,9'd294,9'd311,9'd16,9'd315,9'd299,9'd318,9'd267,9'd318,9'd294,9'd299,9'd269,9'd265,9'd0,9'd260,9'd3,9'd261,9'd268,9'd285,9'd326,9'd19,9'd303,9'd0,9'd81,9'd329,9'd339,9'd328,9'd372,9'd91,9'd39,9'd306,9'd34,9'd30,9'd68,9'd25,9'd277,9'd279,9'd270,9'd282,9'd0,9'd258,9'd260,9'd3,9'd257,9'd262,9'd6,9'd261,9'd71,9'd35,9'd382,9'd267,9'd331,9'd294,9'd300,9'd38,9'd407,9'd375,9'd310,9'd35,9'd316,9'd55,9'd258,9'd298,9'd28,9'd68,9'd10,9'd1,9'd3,9'd264,9'd0,9'd3,9'd1,9'd257,9'd267,9'd258,9'd265,9'd3,9'd313,9'd285,9'd25,9'd8,9'd21,9'd17,9'd18,9'd37,9'd55,9'd266,9'd266,9'd272,9'd9,9'd25,9'd3,9'd7,9'd0,9'd10,9'd1,9'd4,9'd9,9'd6,9'd17,9'd0,9'd6,9'd8,9'd261,9'd0,9'd0,9'd5,9'd265,9'd11,9'd25,9'd0,9'd12,9'd23,9'd24,9'd44,9'd15,9'd8,9'd1,9'd5,9'd9,9'd8,9'd271,9'd12,9'd1,9'd3,9'd14,9'd3})
	) SNN (
		.clk(clk),
		.pixels(pixels),
		.start(start),
		.neuron_out(neuron_out)
	);

	initial begin
		integer i;
		integer j;
		for (j = 0; j < 1038; j = j + 1) begin
			// set pixels
			
        if (j == 0) begin
            pixels = 784'b0000000000000000000000000000000000000010000000000000000000000000011100000000000000000000000011110000000000000000000000001111100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000010000000000000011100000111111100000000000001111111111111110000000000000011111111000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000011111111111000000000000000111100000001100000000000000111000000000011000000000000110000000000001100000000000110000000000000100000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000001100000000000000000000000000011100000000000000000000000000111111111111100000000000000000011111111000000000000000000000111100000000000000000000000111000000000000000000000000111000000000000000000000000111000000000010000000000000011000000001111000000000000001111111111111000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 2) begin
            pixels = 784'b0000000000110000000000000000000000000111100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001110000000000000000000000000011110011000000111000000000001111111111111111110000000000000111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 3) begin
            pixels = 784'b0000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000001000000000000000000000000000100000000000000000000000000111110000000000000000000111111110000000000000000000111000110000000000000000000000000011000000000000000000000000001100000000000000000000000000011000000000000000000000000001110100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 4) begin
            pixels = 784'b0000000000000000000000000000000000000000001000000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000111110000000000000000111111111110000000000000000001111110000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 5) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000111111111010000000000000001111110000011000000000000000111100000001100000000000000011100000000110000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000001111000000000000000000000000011111110000000000000000000000111111111000000000000000000000011111100000000000000000000001111100000000000000000000011111000000000000000000000111110000000000000000000000011100000000000000000000000001110000000001111000000000000111111111111111100000000000001111111111110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 6) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000011111111111000000000000000111111111100000000000000000111111000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001111000110000000000000000000011111111100000000000000000001111111110000000000000000000111111111000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011111110000000000000000000000111111100000000000000000000000111111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 7) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111110000000000000000000000001111111000000000000000000000001111100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000100000000000000000000001110110000000000000000000000011111000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 8) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011101110000000000000000000001111111110000000000000000000011111111100000000000000000000000001110000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 9) begin
            pixels = 784'b0000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000001000000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000111111000000000000000011111111111100000000000000001111111111110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 10) begin
            pixels = 784'b0000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000001110000000000000000000000000111100000000000000000000000001111000000011000000000000000111111111111110000000000000001111111111111000000000000000001111111111000000000000000000011111111100000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 11) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111111000000000000000000011111111100000000000000000011111100111000000000000000011111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000000110000000000000000000000000011110000000000000000000000000111111100000000000000000000000011111100000000000000000000000011110000000000000000000000011111000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001111111111000000000000000000001111111110000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 12) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111111100000000000000000111110000000000000000000000111100000000000000000000000011100000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000001111000001111000000000000000000111111111000000000000000000000111110000000000000000000000011100000000000000000000000011100000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001100000111000000000000000000011111111100000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 13) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000001111111110000000000000000001111001111110000000000000001110000001111100000000000000111000000111110000000000000011100000010000000000000000001110000000000000000000000000111000000000000000000000000001111110000000000000000000000111111100000000000000000000011111110000000000000000000000111100000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011111111100000000000000000000111111110000000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 14) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111111000000000000000000001110011110000000000000000001110000011111000000000000000111000000111100000000000000011100000001110000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111001000000000000000000000011111110000000000000000000000111111000000000000000000000111110000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001100000011110000000000000000110011111111000000000000000011111111000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 15) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111111000000000000000011111101111100000000000000011111111111110000000000000001111111111110000000000000000111110000000000000000000000011100000000000000000000000001110000000000000000000000000011100000000000000000000000001111111110000000000000000000011111111000000000000000000011111000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000110001111000000000000000000011111111000000000000000000000111111000000000000000000000111110000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 16) begin
            pixels = 784'b0000000000000000000000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001100000110000000000000000001110001111100000000000000000110001111100000000000000000111111111100000000000000000011111110000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 17) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000011111111111000000000000000011111100111110000000000000011111100000111000000000000011111111111111100000000000001111111111111110000000000000111000000011110000000000000011100000000000000000000000001110000000000000000000000000111100111000000000000000000001111111110000000000000000000011111111000000000000000000001111111000000000000000000001111000000000000000000000001111000000000000000000000000111111111000000000000000000011111111100000000000000000001111111100000000000000000001111100000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 18) begin
            pixels = 784'b0000000000000000000000000000000000000000000000001000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000011110000000000000000111111111110000000000000000011111111100000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 19) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000111111111110000000000000001111111011111100000000000000111100000001111000000000000111111111111111000000000000011111111111111100000000000001111100110011000000000000000110000000000000000000000000011000000000000000000000000001110000110000000000000000000011110111100000000000000000001111111110000000000000000001111111111000000000000000001111100000000000000000000011110000000000000000000000001110000110000000000000000001110001111100000000000000000111111111111000000000000000001111111111000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 20) begin
            pixels = 784'b0000000000000000000000000000000000000000000000001000000000000000000000000001100000000000000000000000000100000000000000000000000000110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000001111000000000000000111111011111100000000000000011111111110000000000000000001111000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 21) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000001111111100000000000000000011111100000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001111111000000000000000000000111111110000000000000000000111111110000000000000000000111100100000000000000000000111100000000000000000000000011000000000000000000000000001100000000000000000000000000111011100000000000000000000011111110000000000000000000001111110000000000000000000001110000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 22) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000110000000000000000011111111111000000000000000011111111110000000000000000001110000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 23) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000011111110000000000000000001111111111100000000000000001111110001110000000000000001111111000111000000000000000111111111111000000000000000011111111111100000000000000001110000010000000000000000000111000000000000000000000000011111110000000000000000000001111111000000000000000000000111111100000000000000000001111101000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001111111100000000000000000000011111110000000000000000000001111110000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 24) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000011000000000000011100000001111100000000000001111111111111110000000000001111111111100000000000000000111110011100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 25) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000011111111110000000000000000001111111111110000000000000001111000000011100000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000100000000000000000000011111111000000000000000000011111111100000000000000000011111001100000000000000000001100000000000000000000000001110000000000000000000000000111000100000000000000000000011111111000000000000000000001111111000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 26) begin
            pixels = 784'b0000000000000000000000000000000000000000000000100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111011111110000000000000000111111111111000000000000000011111101100000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 27) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000001111111111000000000000000001111000011110000000000000001111000000111100000000000001111111111111110000000000000111111111111111000000000000011100000000110000000000000001110000000000000000000000000111000000000000000000000000001111111000000000000000000000111111100000000000000000000111111110000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011111110000000000000000000000111111100000000000000000000111110000000000000000000000111000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 28) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000100000000000000011100000001111000000000000001111111111111100000000000001111111111111100000000000000111111111110000000000000000011111000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 29) begin
            pixels = 784'b0000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000110000000000000011110000000111100000000000001110000000111110000000000001110000000111110000000000000111000001111110000000000000011111111111100000000000000001111111111000000000000000000011001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 30) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000001000000000000000001100000011110000000000000001111110011110000000000000000111111111110000000000000000111111111100000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 31) begin
            pixels = 784'b0000000000000000000000000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000001000000000000000001110000011110000000000000001110000111111000000000000000111111111111000000000000000011111111100000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 32) begin
            pixels = 784'b0000000000000000000000000000000000000000000001000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000111100000000000000001111111111110000000000000000011111111110000000000000000000011110000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 33) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000010000000000000000001100000111100000000000000001110001111100000000000000000110111111100000000000000000111111110000000000000000000011111000000000000000000000011110000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 34) begin
            pixels = 784'b0000000000000000000000000000000000000000000000100000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000011110000000000000011100001111111000000000000001110001111111000000000000000111111111110000000000000000011111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 35) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000111111111100000000000000000111110000110000000000000000111111111111100000000000000111111111111110000000000000011100000111111000000000000001100000000001000000000000000110000000000000000000000000011100000000000000000000000001111111100000000000000000000111111110000000000000000001111111110000000000000000001111000000000000000000000000110000000000000000000000000011111010000000000000000000011111111000000000000000000001111111000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 36) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111110000000000000001111111111111000000000000000111111101111110000000000000011101111111111000000000000011100000000000000000000000001110000000000000000000000000011100000000000000000000000001111000011110000000000000000011111111111000000000000000001111111111100000000000000000111110000000000000000000000111100000000000000000000000011100000000000000000000000001100000000000000000000000000111100111000000000000000000011111111100000000000000000001111111000000000000000000001111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 37) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000011111111111100000000000000111111011111100000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111111000000000000000000001111111110000000000000000001111111111000000000000000011111000000000000000000000001110000000000000000000000001111000000000000000000000000111011110000000000000000000011111111100000000000000000001111111100000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 38) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111111111110000000000001111110001111111000000000001111100000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000011111111111000000000000000000111111111100000000000000000001111111100000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111000000000000000000000000111000000000000000000000000011111100000000000000000000001111111111111100000000000000011111111111110000000000000000000011101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 39) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000010000000000000000011110000011000000000000000000111110011100000000000000000001111111110000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 40) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000011111111111100000000000000011111100111111000000000000011110000000011100000000000011110000000001110000000000011110000000000011000000000001110000000000000000000000001110000000000000000000000000011000000000000000000000000001110000000000000000000000000111000010000000000000000000001111111100000000000000000000011111110000000000000000000001111100000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011101111110000000000000000001111111110000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 41) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000111000001000000000000000000001100001100000000000000000000011101110000000000000000000000111110000000000000000000000001111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 42) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000011111111000000000000000000111100001111000000000000000111000000011100000000000000011000000000111000000000000011100000000011100000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000000111101110000000000000000000001111111000000000000000000001111111000000000000000000011111000000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000001111111111111000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 43) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000110000000000000001110000000110000000000000000011111000011000000000000000000001111011100000000000000000000001111100000000000000000000000011110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 44) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000011000000000000000011100000011100000000000000001110000001110000000000000000111000011110000000000000000001110001110000000000000000000111111111000000000000000000001111111000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 45) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000001110000000000001111111111111111000000000000011111111111111110000000000000001001111111111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 46) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000100000000000000000001111000111000000000000000000011111011100000000000000000000111111110000000000000000000000111111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 47) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111111110000000000000001111100001111100000000000000111000000000000000000000000011000000000000000000000000001110000000000000000000000000111000000000000000000000000001110000000000000000000000000111110000000000000000000000000111111100000000000000000000001111110000000000000000000001111110000000000000000000001111000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001111111111100000000000000000111111111110000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 48) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001111111000000000000000000001110001110000000000000000001110000001110000000000000000110000000011000000000000000011000000000000000000000000001110000000000000000000000000011000000000000000000000000001110000000000000000000000000011110000000000000000000000000011111110000000000000000000000111111000000000000000000001111100000000000000000000001111000000000000000000000001110000000000000000000000001100000000000000000000000001100000001000000000000000000110000111100000000000000000011111111110000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 49) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000100000000000000001100000000110000000000000000111110000011000000000000000000111111111100000000000000000000011111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 50) begin
            pixels = 784'b0000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000000111111111111100000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 51) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111111100000000000000000111000001111100000000000000011000000001110000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000000111011100000000000000000000011111110000000000000000000001111110000000000000000000011111000000000000000000000001111100100000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000001110000000000000000011110001111100000000000000000111111111100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 52) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111111000000000000000001111000111000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011100000000000000000000000001110000110000000000000000000011111111100000000000000000000111111100000000000000000000111110000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000111111111100000000000000000001111111111000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 53) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111110000000000000000001111000001100000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011100000000000000000000000000111000000000000000000000000001111000100000000000000000000011111110000000000000000000001111111000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 54) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111111110000000000000000011110001111110000000000000111100000000111100000000000011100000000000100000000000001110000000000000000000000000111000000000000000000000000001111000000000000000000000000011111110000000000000000000000111111100000000000000000000111111000000000000000000001111000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000110000000000000000000011111011111000000000000000000111111111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 55) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000001111111111111100000000000011110000000000000000000000011110000000000000000000000001100000000000000000000000000111000000000000000000000000000111110000000000000000000000001111111100000000000000000000111111111000000000000000001111100000000000000000000001111000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111111111100000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 56) begin
            pixels = 784'b0000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000010000000000000000000111111111000000000000000000011111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 57) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001110011111100000000000000001110000001111000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000011000000000000000000000000001111110000000000000000000001111110000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000011100000000000000000000000000111111110000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 58) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000001100000000000000000000000000111100000000000000000000000001111100000000000000000000000001111111000000000000000000000001111111100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 59) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000001111100110000000000000000000001111011000000000000000000000001111100000000000000000000000011100000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 60) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111000100000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000001101000000000000000000000000111110000000000000000000000011110000000000000000000000011100000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000000100000011110000000000000000011001111111000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 61) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000011001111000000000000000000001111111000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 62) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111111100000000000000000001110000011000000000000000001100000000110000000000000001110000000001100000000000000110000000000010000000000000011000000000001000000000000001100000000000000000000000000110000000000000000000000000011111100000000000000000000000111111000000000000000000000111110000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000001110000000000000000000000000011111111100000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 63) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000001100000000000000000001111000110000000000000000000011111111000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 64) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000111111110000000000000000000111111111100000000000000000011110001111000000000000000011110000001110000000000000001110000000011000000000000000110000000000100000000000000011000000000010000000000000001110000000000000000000000000111100000000000000000000000001111100000000000000000000000011111111100000000000000000000111111111000000000000000000011111111100000000000000000011111000000000000000000000011111000000000000000000000001111100000011000000000000000111111111111100000000000000001111111111100000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 65) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000001000000000000000011111111111100000000000000001111111111110000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 66) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000001111111100000000000000000011111111111100000000000000001111100001111000000000000000111100000011100000000000000111100000000110000000000000011110000000011000000000000001111100000001100000000000000011111110000000000000000000000111111100000000000000000000000111111101111100000000000000001111111111110000000000000000001111111110000000000000000001111111110000000000000000001111110000000000000000000001111100000000000000000000000111110000000000000000000000011111111111111000000000000000111111111111000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 67) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111110000000000000000000000111100000000000000000000000111110000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000111100000000111000000000000111110000000011111111100111111111000000001111111111111111111000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 68) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000001111111111000000000000000011111111111110000000000000011111111000111100000000000001111100000001110000000000000111000000000011000000000000011100000000001100000000000001110000000000000000000000000111100000000000000000000000001111000000000000000000000000111111000000000000000000000000111111000000000000000000000001111111111000000000000000001111111111100000000000000001111111000000000000000000001111110000000000000000000000111110000000000000000000000001111111111100000000000000000011111111111100000000000000000001100111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 69) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000011111000000000000000000000011111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111110000000000000000000001111110000000000000000000001111111000000000000000000000111111000000000000000000000111111000000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000011111111111111111100000000001111111111111111110000000000011111111111111111000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 70) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111000000000000000001111111111111000000000000001111000000011100000000000000111100000000011000000000000111100000000001100000000000011100000000000010000000000001110000000000000000000000000111000000000000000000000000001110000000000000000000000000111000111100000000000000000011111111111000000000000000000111111111100000000000000000011111111100000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011111000000000000000000000000111111111110000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 71) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111111000000000000000000000111111000000000000000000000111111000000000000000000000011111000000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000111000000000011111000000011111100000000000111111111111111110000000000011111111111111100000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 72) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000111100000000011100000000011111100000000001111111111111111100000000000111111111111111100000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 73) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000001111000000000001100000000000111111111111111100000000000001111111111111100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 74) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000111000000000000000011110000111100000000000000001111111111111000000000000000001111111111000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 75) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000100000000000001111000000000111100000000000111111111111111100000000000001111111111111100000000000000001111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 76) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111110000000000000000001111111111100000000000000001111000001111000000000000001111000000011000000000000001111000000001100000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001111111110000000000000000000011111111100000000000000000001111111100000000000000000000111111000000000000000000000011100000000000000000000000011100000111110000000000000001111011111111000000000000000011111111110000000000000000001111111111000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 77) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111110000000000000000001111111111110000000000000001111100001111100000000000000111100000001111000000000000111000000000011100000000000011100000000000110000000000001110000000000001000000000000011000000000000000000000000001110000000000000000000000000011100000000000000000000000000111111100000000000000000000001111111100000000000000000000111111110000000000000000000111111110000000000000000000111100000000000000000000000011110000000000000000000000001111110000000000000000000000011111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 78) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000111111000000000000000000001111111111000000000000000000111100011110000000000000000111000000011000000000000000011100000000100000000000000001110000000010000000000000000111000000000000000000000000011110000000000000000000000000111000000000000000000000000001111000000000000000000000000011111100000000000000000000001111111000000000000000000001111111100000000000000000001111100000000000000000000000111000000000000000000000000011100000000000000000000000001111111110000000000000000000011111111000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 79) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001111100000000000000000000000011111111111111100000000000000111111111111110000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 80) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000111111100000000000000000001111111111000000000000000001111100001100000000000000001111000000111000000000000000111000000001100000000000000011100000000110000000000000001110000000001000000000000000011000000000000000000000000000110000000000000000000000000011100000000000000000000000000111111000000000000000000001111111110000000000000000001111111110000000000000000001111000000000000000000000000111000000000000000000000000011110000000000000000000000000111111111110000000000000000001111111111000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 81) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000111111110000000000000000000111111111100000000000000000111000000110000000000000000111000000011000000000000000011100000000100000000000000001110000000000000000000000000111000000000000000000000000001110000000000000000000000000011000000000000000000000000000111000100000000000000000000001111110000000000000000000011111111000000000000000000011111000000000000000000000011110000000000000000000000001110000000000000000000000000111100000000000000000000000001111111000000000000000000000011111110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 82) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000111111110000000000000000001111110111100000000000000001111000000111000000000000000111000000001110000000000000011100000000011000000000000001110000000000100000000000000111000000000000000000000000001110000000000000000000000000111000000000000000000000000001111111000000000000000000000111111110000000000000000000111111111000000000000000001111100111000000000000000000111000000000000000000000000011000000000000000000000000001110000000000000000000000000111100001111000000000000000001111111111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 83) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000011111111000000000000000000011110001110000000000000000011100000011100000000000000011100000000110000000000000001110000000001100000000000000110000000000110000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000000111111100000000000000000000111111111000000000000000000111111111000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000011100000000000000000000000001111111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 84) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111110000000000000000000111111111110000000000000000011100000111000000000000000011100000001100000000000000001110000000000000000000000000111000000000000000000000000001110000000000000000000000000111000000000000000000000000001111111000000000000000000001111111110000000000000000001111111111000000000000000001111001111000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000001111110000000000000000000000011111110000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 85) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000010000000000000000111000000011100000000000000011100000011110000000000000001110000011110000000000000000111000011110000000000000000111111111110000000000000000011111111110000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 86) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000011000000000000111000000000111100000000000011100000000111100000000000011111000111111100000000000000111111111111110000000000000011111111101110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 87) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000011000000000000000011100000011100000000000000001110000001110000000000000000110000001110000000000000000011000011110000000000000000001111111110000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 88) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000001100000000000000001110000001110000000000000000111000000111000000000000000011110001111000000000000000001111111111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 89) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111110000000000000000011111111111100000000000000011110000000110000000000000001111000000011000000000000000111000000000110000000000000111100000000000000000000000011110000000000000000000000000111000000000000000000000000011100000000000000000000000001111100001111100000000000000011111111111110000000000000000011111111111000000000000000000011111110000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001111100111000000000000000000011111111100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 90) begin
            pixels = 784'b0000000000000000000000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011111111111111000000000000001111111111111100000000000000111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 91) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111110000000000000000111111111111100000000000000111110000001111000000000000111100000000001100000000000111100000000000010000000000111000000000000011000000000011100000000000011100000000001100000000111000000000000000110000011111100000000000000011100111111100000000000000000011111111110000000000000000000111111100000000000000000000111100000000000000000000000111100000000000000000000000111000000010000000000000000011000001111100000000000000001100111111100000000000000000011111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 92) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001111111111111110000000000001111111111111111000000000000111111010000011100000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 93) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000001111111110000000000000000011111100011100000000000000111110000000011000000000000111000000000000100000000000111000000000000011000000000111000000000000001100000000011000000000000000010000000001100000111000000001000000000110001111110000000000000000011111111111000000000000000000011111100000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000001110000000000000000111000001111000000000000000011111111111000000000000000000111111111000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 94) begin
            pixels = 784'b0000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000011111100000000000111000111111111110000000000011111111111111111000000000000111111111111111100000000000001100000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 95) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000100000000000000000011100000011000000000000000001100011111110000000000000001111111111111100000000000000111111111111110000000000000001111110011111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 96) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000111110000000000000001110011111111110000000000000111111111111111000000000000011111111100111100000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 97) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111100000000000000000000011111110000000000000000000011111001000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000011110000000000000000000000000111111110000000000000000000001111111100000000000000000000001111110000000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011111111000000000000000000000111111100000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 98) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000001111111111100000000000000011111111111110000000000000011111100000111100000000000011111000000011100000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000000110000011110000000000000000111000111111000000000000000011111111111100000000000000000111111111000000000000000000001111111000000000000000000000111110000000000000000000000111110011000000000000000000011110001100000000000000000011110001110000000000000000011111111111000000000000000001111111111000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 99) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000011110000010000000000000000001111111111111111000000000000111111111111111110000000000001111111111001111000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 100) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000011000000000000001100111111111110000000000000111111111111110000000000000011111111111100000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 101) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000001111111100000000000000000011111111111000000000000000111111000011110000000000000111100000000011100000000000011100000000000111000000000001111100000000000000000000000011111111100000000000000000000011111110000000000000000000000111111000000000000000000000111111000000000000000000000111110000000000000000000000111000000000000000000000000111100011000000000000000000111111111110000000000000000011111111110000000000000000001111111110000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 102) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001111111111000000000000000000111111111100000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 103) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000001111111100000000000000000011111111111000000000000000111111110001110000000000000111110000000011100000000000111110000000000110000000000111110000000000001100000000111100000000000000110000000011100000011000000011000000001110001111110000000000000000111111111111000000000000000001111111111000000000000000000001111110000000000000000000001111110000000000000000000001111100000000000000000000001111100001100000000000000000111100111111000000000000000011111111111000000000000000000111111111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 104) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000001111111110000000000000000011111101111100000000000000011110000000110000000000000011110000000000000000000000011110000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000010000000000000000001111111111100000000000000000001111111110000000000000000000001111110000000000000000000001111110000000000000000000001111100000000000000000000001111000000000000000000000000111000010000000000000000000011111111100000000000000000001111111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 105) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000001110000000000011000000000001111000000000011110000000111111100000000001111111101111111110000000000111111111111100000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 106) begin
            pixels = 784'b0000000000000000000000000000000000000000000100000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011111111111111000000000000000111111111111100000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 107) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111111000000000000000011111111111100000000000000111111000000110000000000000111110000000001100000000000011100000000000010000000000011100000000000000000000000000111101111110000000000000000011111111111000000000000000000111111111000000000000000000001111111000000000000000000001111110000000000000000000001111100000000000000000000001111100000000000000000000001111000000000000000000000001111000011110000000000000000111101111111000000000000000011111111111100000000000000001111111110000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 108) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000110000011111000000000000000111111111111100000000000000011111111100000000000000000011110000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 109) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011111000000000000000000000001111111111111111000000000000111111111111111110000000000001100001111001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 110) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000001111111111100000000000000011111000001111000000000000011110000000001100000000000011100000000000111000000000011100000000000011000000000011100000000000001100000000001100000000000000110000000001100000001111000010000000000010000111111100001100000000001101111111000000100000000000011111110000000000000000000000111100000000000000000000001111000000000000000000000000111000000000000000000000000111100011100000000000000000011111111110000000000000000000111111111000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 111) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000111111111100000000000000000111111111110000000000000000111100001000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000011100000000000000000000000001110000111000000000000000000011111111100000000000000000000111111100000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001100000000000000000000000000111111111100000000000000000011111111110000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 112) begin
            pixels = 784'b0000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000110000000000000000011100000111000000000000000001110000011110000000000000001111000001111000000000000000111000000111100000000000000011111111111110000000000000001111111111110000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 113) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000011111111111100000000000000011111111111110000000000000111110000011100000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000001110000000000000000000000000111000000000000000000000000011111000001100000000000000000111111111110000000000000000000111111110000000000000000000000111110000000000000000000000011110000000000000000000000001110000000110000000000000000111000011111000000000000000011111111111000000000000000001111111110000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 114) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000011000000000000000000000000011100000000000000000000000001110001100000000000000000000110000110000000000000000000111000011000000000000000000011000011100000000000000000011110001110000000000000000001111111110000000000000000000100011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 115) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000001110000000000000000011100000111000000000000000001110000111100000000000000001110000011110000000000000001110000001110000000000000001111000001111000000000000000111111111111000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 116) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000011111111111100000000000000111111111111110000000000000111110000000011000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011111000011110000000000000000111111111111000000000000000000011111111000000000000000000000111111000000000000000000000111110000000000000000000000111110000000000000000000000111100000000000000000000000111110000000010000000000000111110000011111100000000000011111111111111100000000000001111111111111100000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 117) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111111000111000000000000000011111111111100000000000000000011111111110000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 118) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000001111111000000000000000000001111111100000000000000000001111110000000000000000000001111100000000000000000000001111100000000000000000000001111000000000000000000000001111100000000000000000000000111100001110000000000000000011100111111000000000000000001111111111100000000000000000011111111100000000000000000000011111000000000000000000000011111000000000000000000000011111000000000000000000000011111000001000000000000000001111000111110000000000000000111111111110000000000000000011111111100000000000000000000111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 119) begin
            pixels = 784'b0000000000000000000000000000000000000000110000000000000000000000000111100000000000000000000000111110000000000000000000000011111000000000000000000000001111100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000001100000000000000011100000001110000000000000011110000000111000000000000001111000000011100000000000000111111111011110000000000000001111111111111000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 120) begin
            pixels = 784'b0000000000000000000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000011000000000000000111000000001100000000000000011100000001110000000000000001110000000111000000000000001111000000111100000000000000111111111111100000000000000011111111111110000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 121) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111110000000000000000011111111111100000000000000001111100001110000000000000001111000000111000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000011000000000000001110000001111100000000000000011111111111110000000000000000111111111100000000000000000000111111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000011100000000000000111111111111110000000000000011111111111100000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 122) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000011100000000000000001111000001110000000000000000111000001111000000000000000111100001111000000000000000011100000111100000000000000001110000011110000000000000001111111111110000000000000000011111111111000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 123) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111100001110000000000000000011111111111111000000000000001111111111111100000000000000111111111000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 124) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111111000000000000000000011111111100000000000000000111111000010000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000011110000000000000000000000001111111110000000000000000000001111111100000000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000000000000011111000000000000000000000111111111111000000000000000111111111111100000000000000111111111011110000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 125) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000011111000000000000111111111111111100000000000011111111111111100000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 126) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111111100000000000000000011111111110000000000000000011111000011000000000000000011110000011100000000000000001110000010000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001111000000110000000000000000011111001111100000000000000001111111111100000000000000000001111111100000000000000000000001111100000000000000000000001111000000000000000000000001111100000000000000000000001111111111111000000000000011111111111111000000000000001111111111100000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 127) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111100000000000000001111111111111000000000000001111110000001110000000000001111100000000010000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000000111000010000000000000000000011111111100000000000000000000111111110000000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000011111000000000000000000000011111000001100000000000000001111000011111000000000000001111111111111100000000000000111111111111000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 128) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000011111111000000000000000000011111111110000000000000000011111101111000000000000000001111000011100000000000000000111000000100000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011110000000000000000000000000111000000000000000000000000011110000000000000000000000000111111100000000000000000000001111110000000000000000000001111111000000000000000000000111111000000000000000000000011100000110000000000000000001111111111000000000000000000111111111100000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 129) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100011000000000000000000001110001100000000000000000000111001110000000000000000000011100111000000000000000000001110011100000000000000000000111001110000000000000000000001111110000000000000000000000111111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 130) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000011111111110000000000000000111111111111000000000000000111100000001100000000000000011100000000100000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000011100000000000000000000000001110011111000000000000000000011111111100000000000000000001111111100000000000000000000011111110000000000000000000011110000000000000000000000001110000000000000000000000000011100000000000000000000000001111111111000000000000000000011111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 131) begin
            pixels = 784'b0000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000100000000000000011100000000111000000000000001110000000011100000000000000111000000011110000000000000011100000001111000000000000001111000001111100000000000000011110000111100000000000000001111111111100000000000000000011111111100000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 132) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000011111111111000000000000000011111111111110000000000000011110000000111100000000000001110000000001110000000000000111000000000111000000000000011100000000111000000000000001110000000011000000000000000111100000000000000000000000001110000000000000000000000000111100011100000000000000000001111111110000000000000000000011111111000000000000000000001111111000000000000000000001111000000000000000000000000111000000010000000000000000011100000011000000000000000001111111111100000000000000000011111111100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 133) begin
            pixels = 784'b0000000000000000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000001000000000000000001110000001110000000000000000111000001111100000000000000111000000111110000000000000011100000111111000000000000001110000011111100000000000000111000011110000000000000000011111111110000000000000000000111111110000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 134) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000011111111000000000000000000011111111110000000000000000011111111111100000000000000001110000011111000000000000001111000000111100000000000000111000000011110000000000000011100000000110000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111100001100000000000000000001111111111000000000000000000011111111100000000000000000000111111110000000000000000000011111111111000000000000000001111111111110000000000000000111111111110000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 135) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111100000000000000000111111111111000000000000000111100000011100000000000000111000000001110000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000011110011100000000000000000000111111110000000000000000000001111110000000000000000000000111100000000000000000000000111100000000000000000000000011100001000000000000000000001110001110000000000000000000111111111000000000000000000011111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 136) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111111000000000000000111111111111100000000000001111000000011110000000000001111000000001111000000000000111000000000110000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000011110001110000000000000000000111111111100000000000000000001111111100000000000000000000111111000000000000000000000111100000000000000000000000011100000000000000000000000001111001111000000000000000000011111111100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 137) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000111111111100000000000000000111111111111000000000000000111100000111100000000000000011100000000000000000000000001110000000000000000000000000011100000000000000000000000001111000000000000000000000000011110000000000000000000000001111100000000000000000000000011111000000000000000000000000111111111100000000000000000001111111110000000000000000000111111100000000000000000001111111000000000000000000011111100000000000000000000001111100000011000000000000000111111111111100000000000000011111111111110000000000000000111110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 138) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111000000000000000001111111111110000000000000000111000000111100000000000000111000000001110000000000000011100000000001000000000000001110000000000000000000000000011100000000000000000000000001111000000000000000000000000011110000000100000000000000000111110011111000000000000000001111111111000000000000000000001111111000000000000000000000011110000000000000000000000001110000000000000000000000000111000000010000000000000000011100000010000000000000000000111111111000000000000000000011111111000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 139) begin
            pixels = 784'b0000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000001100000000000000011000000000110000000000000001100000000111000000000000001110000000011100000000000000111000000011110000000000000011111100011000000000000000001111111111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 140) begin
            pixels = 784'b0000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000011000000000000000000111000011110000000000000000011100001111000000000000000011110001111000000000000000001111001111100000000000000000011111111110000000000000000001111111110000000000000000000111111100000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 141) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000111111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000100000000000000000000110000111000000000000000000111000011100000000000000000011000011110000000000000000001100001111000000000000000000111011110000000000000000000011111110000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 142) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000001111100000000000000000000000111100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000110000000000000000111000000111000000000000000011000000011100000000000000001100000011110000000000000000111111111100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 143) begin
            pixels = 784'b0000000000000000000000000000000000000001111000000000000000000000000111100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000011100000000000000001100000001110000000000000001110000001111000000000000000110000000111000000000000000111000000111100000000000000011111111111000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 144) begin
            pixels = 784'b0000000000000000000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001110000011000000000000000000111000001100000000000000000111100001110000000000000000011100000111000000000000000001110000011000000000000000000111100011100000000000000000001111111110000000000000000000011111110000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 145) begin
            pixels = 784'b0000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000110000000000000000111000000111100000000000000011100000011110000000000000001100000011111000000000000001111111111111100000000000000111111111110000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 146) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000011111111100000000000000000011111111111100000000000000011110000011110000000000000001110000000111100000000000001110000000001111000000000000111000000000011100000000000001110000000001110000000000000111000000000000000000000000001110000000000000000000000000111100000000000000000000000001111111100000000000000000000111111110000000000000000000011111111000000000000000000011111111000000000000000000001111100000000000000000000000111111111000000000000000000001111111111100000000000000000000111111111000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 147) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000111111100000000000000000000111111111000000000000000000111100111110000000000000000011100000111100000000000000001110000001111000000000000000111000000011110000000000000011100000000111100000000000000111000000001100000000000000001110000000000000000000000000111100000000000000000000000001111100000000000000000000000011111100000000000000000000011111110000000000000000000011111100000000000000000000001111100000000000000000000000011111100011000000000000000000111111111110000000000000000001111111111000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 148) begin
            pixels = 784'b0000000000000000000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000001100000000000000000011100000111000000000000000001100000111100000000000000000110000011110000000000000000011000011111000000000000000001110011110000000000000000000111111110000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 149) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000001111111110000000000000000000111000111100000000000000000111000000111000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000000110000000000000000000000000011000000000000000000000000001110011000000000000000000000011111100000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000001000000000000000000011000000100000000000000000001100000110000000000000000000111001111000000000000000000001111111000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 150) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111110000000000000000011111111111110000000000000001111100011111000000000000001111000000011100000000000000011100000000110000000000000001110000000000000000000000000111000000000000000000000000001110000000000000000000000000111110000000000000000000000001111110000000000000000000000011111110000000000000000000000111111000000000000000000000001111100000000000000000000011111110000000000000000000011111111111000000000000000000111111111111100000000000000001111111111110000000000000000000000001111100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 151) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000011111111000000000000000000011111111111000000000000000011110000011111000000000000001110000000001110000000000000111000000000011000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110001100000000000000000000011101110000000000000000000001111111000000000000000000000111111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111111111111100000000000000111111111111110000000000000011111110001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 152) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100011000000000000000000001110001100000000000000000001110000110000000000000000000111000011100000000000000000011100011110000000000000000001111111110000000000000000000011111111000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 153) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000001110000000000000000011100000111000000000000000001110000011000000000000000000111000011100000000000000000011100001110000000000000000001110000110000000000000000000011100011000000000000000000001111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 154) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000011111111111110000000000000111111100000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000000110000000000000000000000000011000011100000000000000000000110111110000000000000000000011111110000000000000000000001111100000000000000000000000011100000000000000000000000001100000000111000000000000000110000000111100000000000000011000000111100000000000000001100001110000000000000000000110001110000000000000000000011111100000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 155) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000001100000000000000000000000000110000000001000000000000000111000000001100000000000000111111111100110000000000000011110000011111000000000000001110000000111100000000000000000000000001110000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 156) begin
            pixels = 784'b0000000000000001001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000001100011100000000000000000000011111110000000000000000000000111111000000000000000000000011100000000000000000000000011000000000000000000000000001000000000000000000000000001100000011100000000000000000111010111111000000000000000011111111111100000000000000000111111011100000000000000000001101001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 157) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111110000000000000000000111100001100000000000000000011000000110000000000000000001100000011000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000001100000000000000000011000111111000000000000000001111111110000000000000000000001111110000000000000000000000001100000000000000000000000001000000000000000000000000001100000000100000000000000000110000111111100000000000000011111111111000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 158) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110001000000000000000000001111111110000000000000000001111111000000000000000000000111111000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 159) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000011111110000000000000000000111110001000000000000000000111100000100000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000011110000000000000000111100111111000000000000000000111111100000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000110000000000000000111000111111000000000000000011111111111000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 160) begin
            pixels = 784'b0000000000000000000000000000000000000000000001110000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000000011111111111111110000000000011111111111111111100000000001111111111000001110000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 161) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000111111111100000000000000001111111101110000000000000011111110000011000000000000001111000000000100000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001110110000000000000000000000111111000000000000000000000011111100000000000000000000001111000000000000000000000001110000000000000000000000001111000000000000000000000000111000000001100000000000000011100000011110000000000000001110011111111000000000000000111111111100000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 162) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000001111111100000000000000000001111110111000000000000000001111000000100000000000000000111000000010000000000000000111000000001000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000011110000000000000000001111111111000000000000000000111111110000000000000000000001111100000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000111111111100000000000000000000111111111100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 163) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111110000000000000000001111111111100000000000000001110000000110000000000000000110000000001100000000000000010000000000000000000000000001000000000000000000000000000110000000000000000000000000011000000000000000000000000001110111000000000000000000000011111100000000000000000000001111110000000000000000000001111110000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000111100000000000000001111111111110000000000000000011111111111000000000000000000011111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 164) begin
            pixels = 784'b0000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001111100000000000000000000000111111110000000000000000000011111111111100000000000000000111111111111000000000000000000111111111110000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 165) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111110000000000000000000111111111000000000000000000111111001000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000000110000000000000000000000000011111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001111100000000000000000000000011111111000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 166) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001111111111100000000000000000111111111111000000000000000001111111111111000000000000000000000001111100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 167) begin
            pixels = 784'b0000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111001111111000000000000000111111111111110000000000000011111111111111000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 168) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111111000000000000000001111111111100000000000000000111110000010000000000000000111100000000000000000000000011100000000000000000000000001100000000000000000000000000111000000000000000000000000001110000000000000000000000000011111100000000000000000000000111111000000000000000000000011111100000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111111111100000000000000000000011101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 169) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000111100000000000000011111111111111000000000000001111111111000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 170) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111111000000000000000000111111111100000000000000000111110000011000000000000000011100000000100000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100011110000000000000000000011111111000000000000000000000111111100000000000000000000011111100000000000000000000001111100000010000000000000001111100000111100000000000001111000000111110000000000000111100011111000000000000000111111111110000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 171) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111100010000000000000000000111111111111000000000000000001111111111100000000000000000111000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 172) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000111111111111100000000000000111111111111111000000000000011111000000011110000000000001110000000000001000000000000110000000000000110000000000001100000000000000000000000000011000000000000000000000000001111000111000000000000000000001111111110000000000000000000011111111000000000000000000000111111000000000000000000000011110000000000000000000000000111000000111100000000000000011111111111110000000000000000111111110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 173) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000011111111100000000000000000011111111111000000000000000011111110001100000000000000011111000000110000000000000001110000000000000000000000000111000000000000000000000000001100000000000000000000000000011000000000000000000000000000111000000000000000000000000000111111000000000000000000000001111110000000000000000000000111111000000000000000000000111111000000000000000000000111111000000000000000000000111110000000000000000000000011110000000000000000000000001111110110000000000000000000000110011111110000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 174) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101000000000000000000000000100010000000000000000001100000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000000000000000000110000000000000000000000000011100000000000000000000000000111111000000000000000000000011111110000000000000000000011111111000000000000000000011110000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001111000000000000000000000000011111111000000000000000000000000111111000000000000000000000000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 175) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100001000000000000000000001111111110000000000000000001111111111000000000000000001111111100000000000000000000111110000000000000000000000001110000000000000000000000000110000000011000000000000000111000000011100000000000000011100000011100000000000000001100000001110000000000000000110000001111000000000000000011000000111000000000000000001111000111100000000000000000111111111100000000000000000000001111110000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 176) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000111111111111100000000000001111000000011110000000000000110000000000010000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000011110000000000000000001111111111000000000000000000011111000000000000000000000011100000011000000000000000001111111111100000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001100000000000000000000000001000000000000000000000000001000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 177) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011111100000000000000000111111111110000000000000000011111111100000000000000000000111111000000000000000000000000111000000001110000000000000011100000001111000000000000001110000001111000000000000001110000000111100000000000000111000000111100000000000000011100000011100000000000000001111000011100000000000000000011111111110000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 178) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000001111111111111110000000000001111111111111111000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011000000000000000000000000001110000000000000000000000000111000000000000000000000000001110000000000000000000000000111111111111100000000000000000111111111110000000000000000011111111111000000000000000011111000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000011111100000000000000000000000011111111110000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 179) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000111111111100000000000000000111111111110000000000000000001001110000000000000000000000000110000000011000000000000000111000000011100000000000000011000000001110000000000000011100000001110000000000000001110000000111000000000000000111000000111000000000000000011111000111000000000000000000001111011100000000000000000000001111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 180) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000001111111100000000000000000000111111110000000000000000000011111000000000000000000000000011100000000000000000000000011100001100000000000000000001110001110000000000000000001111000111000000000000000000111000011100000000000000000011100001110000000000000000001111000111000000000000000000111111111000000000000000000000001111100000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 181) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000111111111111000000000000000111101001111110000000000000111000000000010000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000000110000000000000000000000000001110001100000000000000000000011111111000000000000000000001111111000000000000000000001111000000000000000000000011110000000000000000000000011110000000000000000000000011100000000000000000000000001110000110000000000000000000011111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 182) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000001110000000000000000000000000010000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000011011110000000000000000000011111111100000000000000000000101110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000110000000000000000111000000111000000000000000011100000111100000000000000001110000011100000000000000000011110011100000000000000000000001111110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 183) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000011111110000000000000000000011111111100000000000000000001111111100000000000000000000001111000000010000000000000000111100000111100000000000000011110000011110000000000000001110000011110000000000000000111000011111000000000000000111100001111000000000000000011110001111000000000000000001111111111100000000000000000011111111100000000000000000000101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 184) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111111111000000000000001111111111101110000000000001110000000111111000000000000110000000000000000000000000011000000000000000000000000000100000000000000000000000000011000000000000000000000000000110000000000000000000000000001111111000000000000000000000011111100000000000000000000001111000000000000000000000011110000000000000000000000111000000000000000000000000011111111100000000000000000000000001111100000000000000000000000000011000000000000000000000000011000000000000000000000000111000000000000000000000101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 185) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000011111111111111100000000000111110000001111110000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011110000000000000000000000000111111111110000000000000000011111111111100000000000000011111111111110000000000000011110000000000000000000000011110000000000000000000000000110000001000000000000000000011000011110000000000000000001111111111000000000000000000011111111000000000000000000000110111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 186) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000011111000100000000000000000011111111111000000000000000011111111111100000000000000001111111111100000000000000000011111100000000000000000000000011110000000011000000000000001110000000001110000000000000111000000000111000000000000011100000000011100000000000000110000000011110000000000000011000000001111000000000000001110000000111100000000000000111000000011110000000000000011100000001111000000000000001111110000111100000000000000011111111111110000000000000000011111111110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 187) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000001111111111100000000000000000110000111110000000000000000110000001111000000000000000010000000000000000000000000001000000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000011000000000000000000000000000111111000000000000000000000001111110000000000000000000001111000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000000110000000000000000000000000011110000000000000000000000000011111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 188) begin
            pixels = 784'b0000000000000000000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000111110000000000000000000000011111000000000000000000000001110000000000000000000000000110000000000000000000000000011000001100000000000000000001100001110000000000000000001110000111000000000000000000110000011000000000000000000011000001100000000000000000001111101110000000000000000000111111110000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 189) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000111111110000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000011110011000000000000000000000011111110000000000000000000001111100000000000000000000001110000000000000000000000011100000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011111111100000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 190) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000001111111100000000000000000001111111100000000000000000000001110000000000000000000000000011000000001000000000000000001100000001100000000000000000110000001100000000000000000110000001110000000000000000011000001110000000000000000001100000110000000000000000000110000110000000000000000000011110110000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 191) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000001111111111100000000000000001110000011111100000000000001110000000011111000000000001100000000001111110000000001110000000000000111000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000000110000000000000000000000000011110000011110000000000000000011111111110000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011000000000000000000000000001111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 192) begin
            pixels = 784'b0000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111100000000000000000000011111111000000000000000000000111111000000000000000000000000110000001100000000000000000011000000110000000000000000001100000111000000000000000000110000011100000000000000000010000001110000000000000000011000001111000000000000000001100000111000000000000000000111111111000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 193) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000011111110000000000000000000011100111000000000000000000011000001100000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000001100000000000000000001111111111000000000000000000011111111000000000000000000011110000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000001100000000000000000000000000011111100000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 194) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000111111110000000000000000000111111111100000000000000000011111111111000000000000000011111011111000000000000000001111000000100000000000000000111000000000000000000000000001110000000000000000000000000111000000000000000000000000001110000000000000000000000000111111000000000000000000000011111100000000000000000000000111110000000000000000000000011111001111000000000000000001111101111100000000000000000111111111110000000000000000011111111110000000000000000000111111110000000000000000000011111110000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 195) begin
            pixels = 784'b0000000000000000000000000000000000000010000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000010000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001111110000000000000000000000111111111000000000000000000001111111110000000000000000000011111111000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 196) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001111111000000000000000000001111111110000000000000000000111111111000000000000000000011100111100000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000011111111000000000000000000000111111110000000000000000000001111111000000000000000000000111111000000000000000000000011111100010000000000000000001111000011110000000000000000011000011111000000000000000001110111111000000000000000000011111110000000000000000000001111100000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 197) begin
            pixels = 784'b0000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000011110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001111111100000000000000000000011111111111000000000000000001111111111110000000000000000111111111111100000000000000000000000111100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 198) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111000000000000000000111111111110000000000000000011111111111100000000000000001111000011110000000000000000111000000011000000000000000001100000000100000000000000000110000000000000000000000000001100000010000000000000000000111001111110000000000000000011111111111000000000000000000111111111111111000000000000001111111111111100000000000000111111101111110000000000000011100111111110000000000000001111111111110000000000000000011111111110000000000000000001111111100000000000000000000111111100000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 199) begin
            pixels = 784'b0000000000000000000000000000000000000111000000000000000000000000011100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000111000000000000000000000000011111111000000000000000000000111111111000000000000000000011111111110000000000000000000011111111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 200) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000011111111000000000000000000001111111110000000000000000000111111111100000000000000000011000011110000000000000000001100000111000000000000000000110000001100000000000000000011000000000000000000000000001110000010000000000000000000011100011100000000000000000001111111110001000000000000000011111111001110000000000000000111111100111000000000000000001111000111100000000000000000111000111100000000000000000011100011100000000000000000001111111110000000000000000000111111110000000000000000000001111110000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 201) begin
            pixels = 784'b0000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011000000000000000000000000001110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001101111111100000000000000000011111111111000000000000000001111111111100000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 202) begin
            pixels = 784'b0000000010000000000000000000000000011000000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111111110000000000000000000001111111111100000000000000000111111111110000000000000000001111111111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 203) begin
            pixels = 784'b0000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000001000000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000001000000000000000000001111111111111000000000000000111011111111100000000000000000101111100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 204) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000001111111000000000000000000000011111110000000000000000000001111111100000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 205) begin
            pixels = 784'b0000000000000000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001110000000000000000000000000111100000000000000000000000011111111100000000000000000000111111111110000000000000000001111111111000000000000000000000011111100000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 206) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000001111111100000000000000000000111111111000000000000000000111111111100000000000000000011000000011000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000000100000000000000000000000000011100000000000000000000000001111111000000000000000000000011111110000000000000000000001111111000010000000000000000001111100011100000000000000000111000011110000000000000000001100001110000000000000000000111111111000000000000000000001111111000000000000000000000111111100000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 207) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000111111110000000000000000000111111111110000000000000000011111111111000000000000000011111000001100000000000000001110000000010000000000000000010000000000000000000000000001000000000000000000000000000110000000000000000000000000011100000000000000000000000000111111000000000000000000000001111100011100000000000000000011110001110000000000000000001111000111000000000000000000111100011100000000000000000011100011110000000000000000000111111111000000000000000000001111111000000000000000000000011111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 208) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111111111100000000000000000011111111111000000000000000000111111111100000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 209) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000001111110000000000000000000001111111110000000000000000000111001111100000000000000000011000001110000000000000000001100000000000000000000000000110000000000000000000000000001000000000000000000000000000110000000000000000000000000001100000000000000000000000000011111000000000000000000000000111110000000000000000000000001111001000000000000000000000111001100000000000000000000011001111000000000000000000001100111000000000000000000000110111100000000000000000000011111100000000000000000000000111110000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 210) begin
            pixels = 784'b0000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011000000000000000000000000001110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000000100000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000001111100000000000000000000000111111110000000000000000000001111111100000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 211) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111111000000000000000001111111111110000000000000000111000000011100000000000000011000000000110000000000000001000000000001000000000000000100000000000000000000000000011000000000000000000000000001110000000000000000000000000011100000000000000000000000000111111000000000000000000000001111110000000000000000000000011110000011100000000000000001110000111111000000000000000110000111111100000000000000011000111111000000000000000001111111100000000000000000000011111000000000000000000000000111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 212) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111110000000000000000001111111111100000000000000000111100001110000000000000000111000000001000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000001100011000000000000000000000111111110000000000000000000011111110000000000000000000001111111000000000000000000000111110001110000000000000000011110011111000000000000000001110011111100000000000000000011011111000000000000000000001111111000000000000000000000011111000000000000000000000001111000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 213) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111110000000000000000000011111111110000000000000000011110000111100000000000000001110000000110000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000011110000000000000000000000000111111100000000000000000000000111110000000000000000000000001111000000011100000000000000111100000011110000000000000011100000011110000000000000001110000011110000000000000000110000011110000000000000000011100011111000000000000000000111111111000000000000000000011111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 214) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000111111100000000000000000000111111111100000000000000000111100001111000000000000000011100000001110000000000000001110000000011000000000000000111000000000100000000000000001110000000000000000000000000011111111000000000000000000000111111110000000000000000000001111111000000000000000000000011111100000000000000000000001110000001000000000000000001110000001110000000000000000111000011111000000000000000011100011111100000000000000000110011111000000000000000000011111111000000000000000000000111111000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 215) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000011111100000000000000000000000111111110000000000000000000000111111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 216) begin
            pixels = 784'b0000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000000111100000000000000000000000011111111100000000000000000000011111111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 217) begin
            pixels = 784'b0000000000000000000000000000000000000100000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000000110000000000000000000000000010000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001100000000000000000000000000111111111100000000000000000001111111111000000000000000000111111111100000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 218) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001111111000000000000000000001111111100000000000000000000110001111000000000000000000010000001110000000000000000001000000011000000000000000001100000001100000000000000000110000000000000000000000000011000000000000000000000000000110000000000000000000000000011000000000000000000000000000111111100000100000000000000011111110001111000000000000000011111001111000000000000000000111000111000000000000000000011000111000000000000000000001101111000000000000000000000111111100000000000000000000011111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 219) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000011111111000000000000000000011111111110000000000000000001100000111110000000000000001100000000111100000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011100000000000000000000000001111000000000000000000000000011111000000000000000000000000111110000000000000000000000001110000000000000000000000001110000000000000000000000000110000001110000000000000000010000001111000000000000000001100011111000000000000000000111111110000000000000000000011111110000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 220) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000001111110000000000000000000011111111000000000000000000111111111100000000000000000111111111111000000000000000011111110011000000000000000001111100000100000000000000000111111111111100000000000000001111111111110000000000000000111111111111000000000000000001111111111100000000000000000011111111000000000000000000001111111000000000000000000000111111100011110000000000000111111111111111100000000000111111111111111110000000000011111111111111110000000000011111111111111110000000000001111111100000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 221) begin
            pixels = 784'b0000000000000000000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000011111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000001111100000000000000000000001111100000000000000000000000111110000000000000000000000111111000011111100000000000011111111111111111000000000011111111111111111100000000001111111111111111110000000000111111111111111110000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 222) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000011111110000000000000000001111111111100000000000000001111111111100000000000000011111111111110000000000000001111111000000000000000000001111100000000000000000000000111100000000000000000000000011110000000100000000000000001111111111111100000000000000111111111111110000000000000011111111111111000000000000000011111111111100000000000000000001111111000000000000000000001111111001110000000000000001111111111111100000000000001111111111111110000000000000111111111111111000000000000011111111110000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 223) begin
            pixels = 784'b0000000000000000000000000000000000000001110000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001110000001111110000000000000111111111111111000000000000111111111111111100000000000011111111111111100000000000001111111110000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 224) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000111111111100000000000000001111111111110000000000000001111111111111000000000000000111111111111100000000000000011111000001100000000000000001111000000000000000000000000111111111100000000000000000011111111111100000000000000001111111111110000000000000000001111111111000000000000000000011111111100000000000000000000111111100000000000000000000111111100000000000000000000111111100011111000000000001111111111111111100000000000111111111111111110000000000111111111111111111000000000001111111111111111100000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 225) begin
            pixels = 784'b0000000000000000000000000000000000000000111000000000000000000000000111110000000000000000000000011111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000000111110000000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000001111111000000011000000000000111111111111111111000000000011111111111111111100000000001111111111111111110000000000111111111111111110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 226) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000001111111111110000000000000001111111111111000000000000001111111111111100000000000001111110000000000000000000000111110000000000000000000000111110000000000000000000000011111100000000000000000000000111111111000000000000000000001111111111000000000000000000011111111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111111000000000000000000001111111111100000000000000001111111111110000000000000000111111111111000000000000000011111111100000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 227) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000001111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111100011111100000000000000111111111111110000000000000011111111111111000000000000001111111111111100000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 228) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111111110000000000000011111111111111000000000000001111111111111000000000000001111110000000000000000000000111110000000000000000000000011110000000000000000000000001111100000000000000000000000111111111111110000000000000011111111111111100000000000000111111111111110000000000000000011111111111000000000000000000001111111000000000000000000001111111000000000000000000001111111000000000000000000000111111000111110000000000000111111111111111000000000000111111111111111100000000000011111111111111100000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 229) begin
            pixels = 784'b0000000000000000000000000000000000000000001111000000000000000000000011111100000000000000000000001111110000000000000000000001111110000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000100000000000111111111111111110000000000011111111111111111000000000011111111111111111100000000001111111111111111110000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 230) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000000000000011111111111000000000000000011111111111100000000000000011111111111000000000000000011111100000000000000000000001111000000000000000000000000111100000000000000000000000011111111111000000000000000001111111111110000000000000000111111111111000000000000000001111111111100000000000000000001111111110000000000000000000001111110000000000000000000011111100000000000000000000001111100000000000000000000011111110111110000000000000001111111111111000000000000001111111111111100000000000000111111111111110000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 231) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000001111111111000000000000000011111111111100000000000000011111111111110000000000000011111110000000000000000000001111100000000000000000000000111100000000000000000000000011111111110000000000000000001111111111100000000000000000011111111110000000000000000000111111110000000000000000000000111111000000000000000000000111111000000000000000000000011111100010000000000000000011111100011000000000000000001111111111110000000000000001111111111111000000000000001111111111111100000000000000111111111111100000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 232) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111100000000000000000000000111100000000000000000000000111110000000001000000000000011110111111111110000000000001111111111111111000000000000111111111111111100000000000011111111100000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 233) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000011111100000000001111100111111111110000000000111111111111111111000000000111111111111111111000000000011111111111100000000000000000111111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 234) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111100000000000000011111111111111110000000001111111111111111111000000000111111111111111111000000000011111111100000000000000000001111100000000000000000000000111111111111000000000000000011111111111100000000000000000111111111110000000000000000000111111110000000000000000000000111111000000000000000000000111110000000000000000000000111111000000000000000000000111111000000000000000000000111111000011110000000000000111111111111111000000000000011111111111111100000000000001111111111111000000000000000111111110000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 235) begin
            pixels = 784'b0000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000011110011111110000000000000001111111111111110000000000001111111111111111000000000000111111111111111100000000000011111100000000100000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 236) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000111110000000000000000000000011110000001100000000000000011111111111110000000000000001111111111111100000000000001111111111111100000000000000111111111111100000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 237) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111111000000000000000111111111111110000000000000011111100011111000000000000011111000000011000000000000001111000000000000000000000001111000000000000000000000000111110000000000000000000000001111111111110000000000000000011111111111000000000000000000111111111100000000000000000000011111110000000000000000000001111110000000000000000000001111110000000000000000000001111110000000000000000000000111110000000000000000000000111111111110000000000000000011111111111100000000000000011111111111110000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 238) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111111111111000000000000000111111111111110000000000000011111111111111000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 239) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000111111111111000000000000000111111111111100000000000000011111110111110000000000000011110000000000000000000000001111000000000000000000000000011110000000000000000000000001111111111110000000000000000011111111111000000000000000000011111111100000000000000000000111111000000000000000000000011111000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111110000011100000000000000111111111111111000000000000111111111111111100000000000011111111111111100000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 240) begin
            pixels = 784'b0000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111100000000000000000000000011110000000000000000000000011111000001011111000000000001111111111111111100000000000111111111111111110000000000011111111111111110000000000011111111111111100000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 241) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111100111110000000000000000111111111111100000000000000111111111111100000000000000001111111111110000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 242) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111111111111110000000000000111111111111111000000000000011111111111111100000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 243) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000111111111111110000000000000111111111111111000000000000111111100111111000000000000111110000000011000000000000011110000000000000000000000001111100000000000000000000000011111111111110000000000000000111111111111100000000000000001111111111110000000000000000000001111110000000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000011111000000000000000000000011111111111000000000000000011111111111100000000000000011111111111110000000000000011111111111110000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 244) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000001111111110000000000000000111111111111000000000000001111111111110000000000000001111111000000000000000000000111110000000000000000000000111110000000000000000000000011111100000000000000000000000111111111000000000000000000001111111111000000000000000000001111111100000000000000000000011111100000000000000000000001111100000000000000000000011111100000000000000000000011111100000000000000000000111111101111000000000000000011111111111110000000000000011111111111111000000000000011111111111111000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 245) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000011111111100000000000000000011111111110000000000000000011110000111000000000000000011110000001100000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011110111100000000000000000000111111111000000000000000000011111111000000000000000000001111111100000000000000000011111111000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100111110000000000000000011111111111000000000000000000111111111000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 246) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111100000011000000000000000111100000011110000000000000111100000111110000000000000011110001111111000000000000001111111111111000000000000000011111111111000000000000000000111111111000000000000000000000001111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 247) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000111111111100000000000000001111110001111000000000000000111100000011110000000000000111100000000111000000000000011100000000011000000000000001110000000000000000000000000110000000000000000000000000011100000000000000000000000001111111111100000000000000000011111111111000000000000000001111111111100000000000000000111111111100000000000000000111111111100000000000000000111100000000000000000000000011100000000000000000000000001111000000000000000000000000011111111000000000000000000000111111110000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 248) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000010000000000000000011100000111000000000000000011100000011100000000000000001110000011110000000000000000111100111110000000000000000011111111110000000000000000000111111111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 249) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000011111110000000000000000000111111111100000000000000000011110001110000000000000000011100000111000000000000000001100000001110000000000000001110000000111000000000000000110000000001000000000000000111000000000000000000000000001100000000000000000000000000111001100000000000000000000011111111000000000000000000001111111100000000000000000001111111100000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001111111111100000000000000000111111111110000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 250) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000011100000011100000000000000001110000011110000000000000001111000011110000000000000000111111111110000000000000000000111111110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 251) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000111111111000000000000000001111000011110000000000000000111000001111100000000000000011000000000110000000000000001100000000011000000000000000110000000000000000000000000111000000000000000000000000001110001100000000000000000000111111110000000000000000000001111111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000011111000000000000000000000001111111111000000000000000000011111111110000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 252) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000111000000000000000011100000111100000000000000011110000111110000000000000001110000011110000000000000001111000111110000000000000000111000111111000000000000000011111111111000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 253) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111111100000000000000001111100001111000000000000000111000000011110000000000000111000000000111000000000000011000000000011100000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000011100000000000000000011111111111000000000000000001111111111000000000000000000011111110000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000011000000000000000000000000001111111110000000000000000000011111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 254) begin
            pixels = 784'b0000000000000000000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000011000000000000000110000000111100000000000000011000000111110000000000000011100000111110000000000000001110001111111000000000000000111111111111000000000000000011111111110000000000000000000111100010000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 255) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000110000000000000011100000001111000000000000001110000001111100000000000001110000011111110000000000000111000111111110000000000000011111111100111000000000000001111111000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 256) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000001110000000000000001110000001111000000000000001111000111111000000000000000011111111111100000000000000000111111111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 257) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000111111111000000000000000000111101111110000000000000000011000011111000000000000000011100000011110000000000000001110000000011000000000000000111000000001100000000000000011100000000000000000000000001110000000000000000000000000011111110000000000000000000001111111000000000000000000001111111100000000000000000000111011110000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000111000000000000000000011111111100000000000000000000111111110000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 258) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000001111111110000000000000000001111111111110000000000000001111000001111000000000000000111000000011100000000000000011000000000110000000000000001100000000011000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111111110000000000000000000011111111000000000000000000011111111100000000000000000011111000000000000000000000011110000000000000000000000001110000000000000000000000000111000001110000000000000000011110011111000000000000000000111111111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 259) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000100000000000000111000000000111000000000000011100000001111100000000000011110000011111100000000000001111111111111100000000000000011111111111110000000000000000011111100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 260) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000011100000000000000000111000001110000000000000000111000011111000000000000000011111111111000000000000000000111111101100000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 261) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000100000000000000011110000000011000000000000001110000000011110000000000001110000000011110000000000000111000000011111000000000000011100000111111000000000000011110001111111000000000000001111111111111000000000000000111111110011100000000000000000111100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 262) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000011111111100000000000000000111111111111000000000000000111111000111110000000000000011110000000111000000000000001110000000011100000000000000111000000000000000000000000011100000000000000000000000001111000000000000000000000000011111001111100000000000000000111111111110000000000000000001111111110000000000000000000111111000000000000000000000011110000000000000000000000001110000010000000000000000001111000001110000000000000000111000000111000000000000000011111111111100000000000000001111111111100000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 263) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000011111111111110000000000000011111111111111100000000000111110000000111110000000000111100000000000111000000000011100000000000001100000000001100000000000000000000000001110000001100000000000000000111000111110000000000000000011111111110000000000000000000011111110000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011111111111100000000000000011111111111111000000000000001110000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 264) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111100000000000000000011111111111000000000000000011110000111110000000000000001110000000111000000000000001110000000001110000000000000111000000000110000000000000011000000000000000000000000001100000000000000000000000000111000000001000000000000000001110001111110000000000000000111111111111000000000000000001111111110000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000011100000011110000000000000001111011111111000000000000000111111111111100000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 265) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000011111111100000000000000000001111111111100000000000000001111000011111000000000000000111000000111110000000000000111000000001111000000000000011100000000011100000000000001110000000000000000000000000111000011110000000000000000011111111111100000000000000000111111111110000000000000000001111111110000000000000000001111110000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011111111110000000000000000001111111111100000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 266) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001111000000000110000000000000111000000000111000000000000011100000001111100000000000001110000001111000000000000001111100111111100000000000000001111111111100000000000000000011111000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 267) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111111111000000000000000011111111111111000000000000011110000011111110000000000001110000000000111110000000000111000000000000111100000000011100000000000000000000000001110000000000000000000000000011100000000000000000000000001110000000000000000000000000111111111100000000000000000001111111110000000000000000000111111111000000000000000000111110000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011111111110000000000000000000111111111100000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 268) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111100000000000000000000000111110000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000011100000000000000001110000011111000000000000001111001111111000000000000000111111111111000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 269) begin
            pixels = 784'b0000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011111000000001110000000000001111111111111111000000000000111111111111111100000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 270) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000001111110000000000000000000011111110000000000000000000011111100000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111100000000000000000000000001111000110000000000000000000011111111100000000000000000001111111110000000000000000001111111000000000000000000001111100000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001111111111100000000000000000011111111110000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 271) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011110000000000000000000000000111000000000000000000000000011110000001110000000000000000111111111111000000000000000011111111111100000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 272) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111111100000000000000000111111111110000000000000000111111100000000000000000000011100000000000000000000000001100000000000000000000000000011000000000000000000000000001110000000000000000000000000011111111000000000000000000000111111110000000000000000000001111111000000000000000000001111111100000000000000000001111100000000000000000000000111100000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000001111111000000000000000000000011111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 273) begin
            pixels = 784'b0000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000011111000111100000000000000001111111111111110000000000000011111111111111000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 274) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000011111111110000000000000000111111111111100000000000000111111111111110000000000000111111000000110000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000000011110000000000000000000000001111111111100000000000000000011111111110000000000000000000011111111000000000000000000001111111000000000000000000000111100000000000000000000000111100000000000000000000000001100000000000000000000000000111111000000000000000000000011111100000000000000000000000111110000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 275) begin
            pixels = 784'b0000000000001100000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011110000001101110000000000000111111111111111000000000000011111111111111100000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 276) begin
            pixels = 784'b0000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000100000000000100000000000000010000111111110000000000000011111111111111000000000000001111001001111000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 277) begin
            pixels = 784'b0000000000000000000000000000000000000001111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000001111100000000000000111111111111110000000000000011111111111110000000000000001111111111010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 278) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000111111111111000000000000001111111111111110000000000001111111111111111100000000000111111101110011110000000000111100000000000000000000000001100000000000000000000000000111000000000000000000000000011111100011110000000000000000111111111111000000000000000001111111111100000000000000000001111111100000000000000000000111111100000000000000000000011000000000000000000000000001100000000000000000000000000110000000111000000000000000011100011111100000000000000001111111111110000000000000000011111111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 279) begin
            pixels = 784'b0000000000000000000000000000000000000011000000000000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000011100000000000001111111110001110000000000000111111111110111000000000000011110001111111100000000000000000000000111110000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 280) begin
            pixels = 784'b0000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000011100000000000001100000000001110000000000000111000000001111100000000000011111011111111111000000000001111111111111111110000000000111111111111111111000000000001000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 281) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000001110000000000000001111111111111000000000000000100111111111100000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 282) begin
            pixels = 784'b0000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000001110000000000001110000000000111000000000000111000000000111000000000000011111100111111100000000000001111111111111110000000000000111111111111111000000000000001000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 283) begin
            pixels = 784'b0000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000001000000000000011111011100001110000000000001111111111111111000000000000111111111111111100000000000001000110001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 284) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000111111111000000000000000001111111111100000000000000011111111000000000000000000001111000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011111111110000000000000000000111111111000000000000000000000111111000000000000000000000111111000000000000000000000011111000000000000000000000001110000000000000000000000001100000000000000000000000000110000000100000000000000000011111111110000000000000000001111111111000000000000000000011111110000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 285) begin
            pixels = 784'b0000000000000010000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000010000000000000000000000000011000000000001000000000000001100000000011100000000000000111111111111110000000000000011111111111111000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 286) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111000000000000000000111111111110000000000000000011111111111100000000000000011111000111110000000000000000110000000001100000000000000011110000000100000000000000000111111110000000000000000000011111111100000000000000000000111111100000000000000000000001111100000000000000000000000010110000000000000000000000001110000000000000000000000001100000000000000000000000000111000000000000000000000000011100000111000000000000000000111110111110000000000000000011111111110000000000000000000111111111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 287) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111110000000000000000001111111111000000000000000000111111111110000000000000000011100000000000000000000000001110000000000000000000000000011110000000000000000000000001111100000000000000000000000011111111110000000000000000000011111111000000000000000000000111111100000000000000000000111111110000000000000000000111110000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000011111111111100000000000000001111111111110000000000000000001111111110000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 288) begin
            pixels = 784'b0000000000000000000000000000000000000000010000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000010000000000000000001100000011000000000000000000110000001100000000000000000011000000010000000000000000001111111111000000000000000000111111111100000000000000000011110000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 289) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000111111100000000000000000000111111110000000000000000000011111100000000000000000000001110000000000000000000000000110000000000000000000000000011100000000000000000000000001111000000000000000000000000011111111100000000000000000000111111110000000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000011000000000000000000000000001100000100000000000000000000111111111000000000000000000001111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 290) begin
            pixels = 784'b0000000000000000000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000110000000000000011100000000011000000000000001110000000001100000000000000111111000001110000000000000001111111111110000000000000000011111111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 291) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000001111111110000000000000000001111111111000000000000000001111111111000000000000000000111110001100000000000000000111100000000000000000000000001100000000000000000000000000111000000000000000000000000001111111000000000000000000000111111100000000000000000000001111110000000000000000000000011111000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000111000111100000000000000000011111111110000000000000000000111111110000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 292) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000111111111100000000000000011111111110000000000000000001111111100000000000000000001111100000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001111000000000000000000000000011111111000000000000000000000111111100000000000000000000001111110000000000000000000001111110000000000000000000000111100000000000000000000000111000000000000000000000000011000000000000000000000000000111000000111000000000000000011111111111100000000000000000111111111110000000000000000000111010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 293) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000111111111110000000000000001111111111111000000000000001111111100111100000000000000111111000000100000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000001111100000111110000000000000011111111111111000000000000000111111111111100000000000000001111111111110000000000000000111111111110000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000000011100001111100000000000000001111111111110000000000000000111111111111000000000000000000011001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 294) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111110000000000000001111111111111100000000000001111111000001110000000000001111100000000001000000000000111100000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000001111000000000000000000000000011111100000000000000000000000111111000000000000000000000011111000000000000000000000011111100000000000000000000001110000000000000000000000000111000000000000000000000000001100000000000000000000000000111111111110000000000000000001111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 295) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000001111111110000000000000000001111111111000000000000000000111111111110000000000000000011111111111000000000000000001100000001100000000000000000111000000010000000000000000011111100000000000000000000000111111000000000000000000000001111100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000011100000000000000000000000001111001100000000000000000000011111111000000000000000000001111111100000000000000000000001111110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 296) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000111111111111000000000000000011111001111110000000000000001110000000010000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100111100000000000000000001111111111000000000000000000111111111000000000000000000011111110000000000000000000001111000000000000000000000001111000000111000000000000001111000000111100000000000000111100011111110000000000000011100111111000000000000000001111111110000000000000000000111111110000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 297) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000001110000000000000000111000001110000000000000000011100001111000000000000000011100001111000000000000000001110000111100000000000000000111100111100000000000000000111111111100000000000000000111100111110000000000000000011100000100000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 298) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111111100000000000000000111111111111100000000000000111100111111110000000000000011100000000111000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001100001100000000000000000000111101111000000000000000000001111111000000000000000000000111111100000000000000000000111100000000000000000000000011110000000000000000000000011100000000000000000000000001110000001000000000000000001111011111100000000000000000111111111110000000000000000011111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 299) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000100000000000000001110000000111000000000000000111000000111100000000000000111000000111100000000000000011100000111100000000000000011111111111100000000000000001111111111100000000000000000111111111000000000000000000111000111000000000000000000011100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 300) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000011111111111110000000000000011100111111111000000000000001110000000011100000000000001110000000000100000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000001111111111100000000000000000011111111110000000000000000000111111110000000000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000111000000000000000011111111111100000000000000001111111111000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 301) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000110000000000000000011000000111000000000000000011100000011100000000000000001100000011100000000000000001110000011100000000000000000111111111110000000000000000111111111110000000000000000011110001110000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 302) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000110000000000000001100000000111000000000000001110000000011100000000000000111000000011100000000000000011001111011100000000000000011111111111100000000000000001111111111110000000000000001111100000110000000000000000111100000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 303) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000111111110000000000000000000111111111100000000000000000111111111111000000000000000011111100011100000000000000001110000000010000000000000000110000000000000000000000000011000000000000000000000000001100000110000000000000000000111001111000000000000000000011111111000000000000000000000111110000000000000000000000011100000000000000000000000011100000000000000000000000011100001100000000000000000001110001111000000000000000000110011111000000000000000000111111110000000000000000000011111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 304) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111000000000000000001111111111110000000000000001111111111111000000000000000111111100111100000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001110001111110000000000000000011111111111000000000000000000111111111000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111001111000000000000000000011111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 305) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000001110000000000000000011000001111000000000000000011100001111000000000000000011100001111000000000000000001110001110000000000000000001111000110000000000000000000111111111000000000000000000111111111000000000000000000011110000100000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 306) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000011111111111110000000000000011111111111111100000000000011111111111111110000000000011111111111111111000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000011110000000000000000000000000111111111110000000000000000001111111111000000000000000000011111111000000000000000000011111000000000000000000000011110000000000000000000000011110000000011000000000000001111111111111110000000000000011111111111111000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 307) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001100000011000000000000000001110000111100000000000000000110000111100000000000000000111000111100000000000000000011111111000000000000000000011111111000000000000000000001110010000000000000000000001110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 308) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000011111111111111000000000000011111100001111100000000000011111000000011100000000000001110000000000100000000000000110000000000000000000000000111000000000000000000000000011100000000001000000000000001110000000111110000000000000011100011111111000000000000000111111111111000000000000000001111111110000000000000000000111100000000000000000000000111100000000000000000000000111100000010000000000000000011100000000000000000000000001110000111110000000000000000111000111110000000000000000001111111100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 309) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000110000000000000000111000000111000000000000000111000000111100000000000000011100001111100000000000000011110000111110000000000000011111110011110000000000000001111111111100000000000000000111001111110000000000000000111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 310) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111111100000000000000001111111111111000000000000001111111111111100000000000001111000011111110000000000000111100000011110000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001100000111110000000000000000111111111111000000000000000001111111111100000000000000000011111111000000000000000000011110000000000000000000000011110000000000000000000000001110000111000000000000000001111011111100000000000000000111111111100000000000000000001111110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 311) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111000000000000000000111111111110000000000000001111111111111000000000000000111111111111100000000000000111100000001110000000000000011100000000000000000000000001110000000000000000000000000111100000111000000000000000011110001111110000000000000000111111111111000000000000000001111111111100000000000000000111111111000000000000000000011110000000000000000000000011110000000000000000000000001110000001000000000000000000111000111110000000000000000011111111110000000000000000001111111110000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 312) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000100000000000000000111000000111000000000000000011100000111100000000000000011100000111100000000000000001111000011100000000000000001111111111100000000000000000111111111100000000000000000111100111100000000000000000011100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 313) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000001111111111100000000000000001111111111111000000000000000111000000001000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011100011100000000000000000001111111110000000000000000000011111110000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000110000000000000000111000001111000000000000000011100011111000000000000000001111111111000000000000000000111111100000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 314) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000001111111111110000000000000001111111111111100000000000001111000111111110000000000011110000000011111000000000001110000000000011100000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000010000000000000000001111000111110000000000000000111111111110000000000000000000111111111100000000000000000011111111000000000000000000011110000111100000000000000001110000111111000000000000001110011111111000000000000000111111111111000000000000000011111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 315) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000001111111111110000000000000000111111111111100000000000000111111111111110000000000000111000000001111000000000000011100000000001000000000000001110000000000000000000000001110000000000000000000000000011000000000000000000000000001110000000000000000000000000111000001110000000000000000011111111111000000000000000000111111111100000000000000000001111111000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001111111100000000000000000000111111110000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 316) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000001110000000000000000000000011100000000000000000000000111100000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000001100000000000000000000000001110000000000000000000000000011100000000000000000000000001111111100000000000000000000001111110000000000000000000001111000000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000011111000011000000000000000001111111111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 317) begin
            pixels = 784'b0000000000000000010000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001111111111111000000000000000111111111111110000000000000011111111111111000000000000000111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 318) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000000000000000000001111000000000000000000000000110000000000000000000000000110000000000000000000000001111000000000000000000000001111000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000110000000000000000111111111111000000000000000001111111111000000000000000000011111100000000000000000000001111000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000001110000000000000000110000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 319) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111110000000000000000001110000001000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000001000000000000000000000000001110000000000000000000000000011111111000000000000000000000011111100000000000000000000001110000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000000110001100000000000000000000011111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 320) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000100000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000001000000000000000000000000001100000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000110101100000000000000000000011111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 321) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000001111100000000000000000000011000000000000000000000000011000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000001100000000000000000001111111110000000000000000000001111100000000000000000000000110000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000000110000000000000000000000000000110000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 322) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001100000000000000000000000011000000000000000000000000111000000000000000000000000110000000000000000000000000110000000000000000000000000010000000000000000000000000011000000000000000000000000001100000000000000000000000000100000000000000000000000000011000000000000000000000000000110000000000000000000000000001111100000000000000000000000111110000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000000100000000000000000000000000000010000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 323) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000000000011000000000000000000000001111100000000000000000000000111100000000000000000000000110000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000001011000000000000000000000000111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 324) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000001000000000000000000000000011000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000011100110000000000000000000000111111000000000000000000000001111100000000000000000000000111100000000000000000000000000000000000000000000000000001000000000000000000000000001100000000000000000000000000011110000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 325) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001000000000000000000000000010000000000000000000000000110000000000000000000000000110000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000000110000011000000000000000000010011111100000000000000000000000111100000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000001100100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 326) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001000000000000000000000000001000000000000000000000000000100000000000000000000000000010000000000000000000000000010000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 327) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110110000000000000000111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 328) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000010100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001111111111000000000000000000111111111100000000000000000001000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 329) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000111100000000000000000000000111110000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000000111000000000000000000000000011100000000000000000000000001111011111000000000000000000011111111110000000000000000000011111110000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 330) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000001000000000000000000000000000000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000011000000000000000000000000000100000110000000000000000000001111111000000000000000000000011111100000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000000110000000000000000000000000001110110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 331) begin
            pixels = 784'b0000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000100000000000000000000000001010000000000000000000000000101000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111000011000000000000000000111110111100000000000000000011111111000000000000000000001110000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 332) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001000000000000000000000000001000000000000000000000000001100000000000000000000000000000000000000000000000000000110000000000110000000000000011000000000111100000000000001100000111111100000000000001110011111111100000000000000111111111111100000000000000001111100001100000000000000000100000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 333) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000100000000000000000000000000110000000000000000000000000110000001100000000000000000010001111010000000000000000011011110000000000000000000001111100000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 334) begin
            pixels = 784'b0000000000000000000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000001110000000000000000000000001111000000000010000000000000111000000000111100000000000011100000000111100000000000001110000000111110000000000000111000000011110000000000000011100000011110000000000000001110000111110000000000000000111111111110000000000000000011111111100000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 335) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000111111100000000000000000000111100011000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000001100000000000000000000000000011010011110000000000000000000001111111000000000000000000000001111000000000000000000000001100000000000000000000000011100000000000000000000000011000000000000000000000000011100000000000000000000000001111111000000000000000000000011111100000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 336) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000011111111000000000000000000111100000111000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000010000000000000011000000000111000000000000011100000000111100000000000011100000000111000000000000001110000001111000000000000000111000011111000000000000000001111111111000000000000000000111111110000000000000000000000000111000000000000000000000000111000011100000000000000000011111111110000000000000000001101111100000000000000000000111111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 337) begin
            pixels = 784'b0000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000100000000000011000000000001110000000000001100000001111111000000000000111111111111111000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 338) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111110000000000000001111000000001100000000000001110000000000011000000000001110000000000001100000000001100000000000000110000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000110000000000000000110000111111000000000000000001111111110000000000000000000001111100000000000000000000000001100000000100000000000000001110000001110000000000000001110000111110000000000000000111111111100000000000000000111111111000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 339) begin
            pixels = 784'b0000000000000000000000000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000111000000011110000000000000011111111111111000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 340) begin
            pixels = 784'b0000000000000000000000000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000011111100000000000011100111111111110000000000001111111111100000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 341) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001110000000000000000000000011110000000000000000000000011100000000000000000000000111100000000000000000000000111100000000000000000000000111000000000000000000000001111000000000000000000000001111000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000000110000000000000000100000000011110000000000000010000000000111111111000011110000000000000001111111111110000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 342) begin
            pixels = 784'b0000000000000000000000000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000000110000000111110000000000000011111111111111100000000000000111111111000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 343) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000011111111111100000000000001111100000000111000000000001111000000000000110000000001110000000000000011000000001110000000000000000000000000111000000000111100000000000001111100011111110000000000000011111111111000000000000000000001111100000000000000000000000111000000000000000000000000111000000000000000000000000111000011111000000000000000011111111111100000000000000011111111111110000000000000000111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 344) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000001111111000000000000000000011111101100000000000000000111110000000000000000000000111100000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000000111100000111111000000000000011111111111111100000000000000011111111110000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011000000000000000000000000001111111111111110000000000000111111111111111000000000000000111111111110000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 345) begin
            pixels = 784'b0000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000001100000000000111000000000001110000000000011000000001111100000000000011111111111111100000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 346) begin
            pixels = 784'b0000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000011100000000000111000000000111100000000000011100011111111100000000000011111111111111000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 347) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000011111111111110000000000001111111000000001100000000001111000000000000010000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000011100000000000000000000000001111000000000000110000000000001111111000111111000000000000001111111111111100000000000000000011111100000000000000000000011100000000000000000000000111100000000000000000000000011000000000000000000000000001100100000000000000000000000111111111111111000000000000000111111111111100000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 348) begin
            pixels = 784'b0000000000000000000000000000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000011111111111001000000000000001111111111111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 349) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111111100000000000000011110000000011100000000000011100000000000110000000000001100000000000000100000000001100000000000000001000000001100000000111000000000000000110000000111100000000000000011000001111100000000000000001110001111000000000000000000011111100000000000000000000000011100000000000000000000000001100000000000000000000000000110000011000000000000000000110000111100000000000000000001111111000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 350) begin
            pixels = 784'b0000000000000000000000000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000010000000000000011000000000011000000000000001100000000111100000000000000111111111111000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 351) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000011111111111111000000000000111110000000000000000000001111000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000011000000000000111100000011111110000000000000111111111111110000000000000000111111000000000000000000000111110000000000000000000000111100000000000000000000000111000000001110000000000000011000000011111100000000000001110000111111111000000000000111111111111100000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 352) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000011110000000000000011000001111110000000000000001111111111100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 353) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000001111111000000000000000000011111111100000000000000000011111111110000000000000000111111100011100000000000000011111000001100000000000000011111000000000000000000000001111100000000000000000000000111101111100000000000000000011111111111000000000000000001111111111000000000000000000111111111000000000000000000011111111000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000000111111111110000000000000000011111111111110000000000000000111111111111000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 354) begin
            pixels = 784'b0000000000000000000000000000000000000000000000111000000000000000000000000111110000000000000000000000111111000000000000000000001111111000000000000000000000001111000000000000000000000001111000000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000000111100000000000000000000001111100000000000000000000000111110000000000000000000000111110000011100000000000000111110001111110000000000000111111111111111000000000000011111111111110000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 355) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000001111111110000000000000000001111110001000000000000000111111000000000000000000000011110000000000000000000000111110000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001111100111000000000000000000111111111100000000000000000000111111110000000000000000001111111000000000000000000001111110000000000000000000000111100000000000000000000000011111000000000000000000000000111111111100000000000000000001111111111000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 356) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000011111111111111000000000000111111111111111110000000000011111111000001111000000000001111110000000001100000000001111000000000000000000000000111110000000000000000000000011111111111000000000000000001111111111100000000000000000111111111110000000000000000111111111100000000000000000111111111000000000000000000011111111110000000000000000000011111111111000000000000000000111111111100000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 357) begin
            pixels = 784'b0000000000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000011111000000000000000000000111111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000001111100000000000000000000001111100000000000000000000001111110000011000000000000001111110000111110000000000001111110000111111000000000001111111001111111000000000001111111111111111000000000000111111111111111000000000000011111111111110000000000000001111000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 358) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000011111111111000000000000000111111111111100000000000000011111000000110000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001111000000110000000000000000111111111111000000000000000001111111111100000000000000000011111111110000000000000000001111111100000000000000000001111111000000000000000000001111110000000000000000000000111110000000000000000000000011111000011111000000000000001111111111111110000000000000011111111111110000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 359) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000000111110000000000000000000000111100001111000000000000000111110001111100000000000000111110111111100000000000000111111111111100000000000000111111111111100000000000000111111111011000000000000000011110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 360) begin
            pixels = 784'b0000000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011110000001110000000000000001110000011111000000000000001111111111111000000000000000111111111100000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 361) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000011111111111100000000000000111111100000111000000000000111110000000011100000000000011110000000000100000000000011110000000000110000000000001110000000000000000000000000111000000000000000000000000011110000000000000000000000000111111000000000000000000000001111111000000000000000000000111111100000000000000000011111111100000000000000000011111110000000000000000000011111100000000000000000000000111111110000000000000000000011111111111100000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 362) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111000000000000000000001111111110000000000000000111111111110000000000000001111111100000000000000000001111110000000000000000000001111100000000000000000000000111000011000000000000000000011111111100000000000000000001111111111000000000000000000111111111000000000000000001111111100000000000000000001111110000000000000000000001111100000000000000000000000111110000000000000000000000011111111100000000000000000000111111111111000000000000000000111111111100000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 363) begin
            pixels = 784'b0000000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000000111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100001110000000000000001111100001111000000000000011111110011111110000000000001111111111111110000000000001111111111111100000000000001111111111111000000000000000111111111010000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 364) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111111000000000000000111111111111110000000000000111111000001111000000000000011111000000001100000000000011111000000001100000000000001111000000000100000000000000111000000000000000000000000111100000000000000000000000001111000000000000000000000000011111111110000000000000000001111111111100000000000000000011111111100000000000000000011111111000000000000000000111111110000000000000000000011111111100000000000000000001111111111000000000000000000111111111000000000000000000001111111110000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 365) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111000000000000000000000000111000000000000000000000000111101111110000000000000000111111111111000000000000000111111111111000000000000000011111011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 366) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000001111110000000000000000000001111110000000000000000000001111111000000000000000000001111111000000000000000000001111110000000000000000000001111110000000000000000000001111110000000000000000000001111110000000000000000000001111110000000000000000000001111110000000000000000000001111110000000000000000000000111110000000000000000000000111111000000000000000000000111111000001110000000000000011111111111111100000000000001111111111111110000000000000111111111111110000000000000001000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 367) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000111111111111111100000000000011111000000001110000000000001110000000000010000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111001110000000000000000000011111111000000000000000000011111111100000000000000000111111100000000000000000000011111000000000000000000000011111000000000000000000000001111111111100000000000000000001111111110000000000000000000000011111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 368) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000001111111100000000000000001111111111110000000000000111111111100000000000000000111111110000000000000000000111111000000000000000000000111110000000000000000000000111110000000000000000000000011110000001110000000000000000111000011111100000000000000001111111111110000000000000000111111111100000000000000000001111111000000000000000000011111110000000000000000000011111100000000000000000000001111100000000000000000000001111111100000000000000000000111111111111110000000000000001111111111111000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 369) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000011111000000000000000000000011111000000000000000000000011111000000000000000000000011110000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000011110000000000000000000000011111000011100000000000000011111111111110000000000000001111111111111000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 370) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111111110000000000001111111100000011000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100011000000000000000000000111111100000000000000000000011111110000000000000000000011111100000000000000000000111110000000000000000000000011100000000000000000000000001111000000000000000000000000111111100000000000000000000000111111100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 371) begin
            pixels = 784'b0000000000000000000000000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000000111100000000000000000000000011110000000000000000000000111100001110000000000000000011100001111100000000000000011100011111100000000000000011111011111110000000000000111111111111000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 372) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110111100000000000011111111111111110000000000111111111111111100000000000011111111110000000000000000011111100000000000000000000001111000000000000000000000000111100000000000000000000000011111000011110000000000000000111111111111000000000000000001111111111100000000000000000111111111100000000000000000111111110000000000000000000111111100000000000000000000111111100000000000000000000011111111111110000000000000001111111111111111110000000000000111111111111111100000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 373) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111110000000000000000001111111111100000000000000001111000111111000000000000000111000000111000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000011111111110000000000000000000011111111000000000000000000000001111000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000000111000010000000000000000000011111111100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 374) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001100000000110000000000000000110000011111000000000000000011111111111000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 375) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111100000000000000000001111110000000000000000000001111000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000001111000000000000000000000000011111111100000000000000000000111111100000000000000000000000111100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000111111000000000000000000000001111110000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 376) begin
            pixels = 784'b0000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000011111111100000000000011111111111111110000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 377) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111111110000000000000001111111111111000000000000001110000000001100000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000000111000111100000000000000000001111111110000000000000000000011111110000000000000000000000111110000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000010000000000000000000111000111000000000000000000001111111000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 378) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000011110000000000000011111111111111000000000000001111111111110000000000000000111110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 379) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000111000000000000000110000000001110000000000000001100000000111000000000000000111111111111100000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 380) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000111100000000000000011000001111110000000000000001111111111110000000000000000111111111100000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 381) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000011111111111000000000000000011111111111100000000000000001111100000100000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001110000000000000000000000000011111111111000000000000000000011111111100000000000000000000111110000000000000000000000001110000000000000000000000000110000000000000000000000000011100000000000000000000000001110001100000000000000000000011111110000000000000000000000111111000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 382) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000001110000000000000001111000111111000000000000000011111111110000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 383) begin
            pixels = 784'b0000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000110000000000000000001100011111000000000000000000111111111100000000000000000011111111000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 384) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001111111111110000000000000000111111111111000000000000000001111111111100000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 385) begin
            pixels = 784'b0000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000001100000000000011100000000000110000000000001110000000000111000000000000111001111000011000000000000011111111111111100000000000001111111111111110000000000000011111111111111100000000000000100000000011100000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 386) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000001100000000000000000011000000110000000000000000001111111111100000000000000000011111111100000000000000000000001110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 387) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000001111111110000000000000000001111111111100000000000000001111110000110000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000011111000110000000000000000000111111111100000000000000000000111111100000000000000000000001111000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111000010000000000000000000011111111000000000000000000000111111100000000000000000000001111110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 388) begin
            pixels = 784'b0000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011110100000000000000000000001111111100011100000000000000111111111111110000000000000011111111111111000000000000001111001111111100000000000000010000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 389) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111110000000000000000001111100111100000000000000000110000000010000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000001100000000000000000000000000111001111000000000000000000001111111000000000000000000000011111100000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011100000000000000000000000000111101100000000000000000000011111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 390) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000011111111110000000000000000011111100111000000000000000011110000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011100000000000000000000000001111000000000000000000000000001111111000000000000000000000011111100000000000000000000000111000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011100000000000000000000000001111111000000000000000000000011111100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 391) begin
            pixels = 784'b0000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000100000000000000001100000000111000000000000000111111111111100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 392) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000111111110000000000000000001111111111000000000000000001111100001000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011100001110000000000000000000111111111000000000000000000001111111000000000000000000000011111000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011000010000000000000000000001111111000000000000000000000011111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 393) begin
            pixels = 784'b0000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000001000000000000000001110000001110000000000000000111111111111000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 394) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111111100000000000000001111111111100000000000000001111110000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011110011110000000000000000000111111110000000000000000000001111111000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111011111000000000000000000011111111110000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 395) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000001111111111110000000000000001111111111110000000000000001111000000000000000000000000111100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111000111000000000000000000011111111000000000000000000000111111100000000000000000000001111100000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001110011100000000000000000000011111111000000000000000000000111111000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 396) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111100000000000000000000111111010000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011000000000000000000000000001111110000000000000000000000011111000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000001101111000000000000000000000111111100000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 397) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111111100000000000000001111111111000000000000000001111000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000001110000000000000000000000000111111100000000000000000000001111110000000000000000000001111110000000000000000000001111000000000000000000000000110000000000000000000000000010000000000000000000000000001111100111000000000000000000111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 398) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111110000000000000000001111111111000000000000000001110000001100000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000110000000000000000000011111111000000000000000000000111111000000000000000000000001111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001111111100000000000000000000111111110000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 399) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000111111000000000000000000001111111110000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000110000000000000000000000000011000000000000000000000000011100001111000000000000000000111111111100000000000000000001111111100000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001111000000000000000000000000001111110000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 400) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000111000000000000000011100000111100000000000000001111000111110000000000000000111111111110000000000000000001111111111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 401) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000111111111000000000000000000111111111100000000000000000111111111110000000000000000111100000000000000000000000111000000000000000000000000011000000000000000000000000011100000010000000000000000000110001111000000000000000000011111111100000000000000000001111111110000000000000000000111111110000000000000000000011111000000000000000000000001110000000000000000000000000110000000000000000000000000011100000000000000000000000001111100000000000000000000000111110000000000000000000000001111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 402) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000011000000000000001110000000011000000000000000111000000011100000000000000011100000001100000000000000001111110001110000000000000000111111111110000000000000000011111111111000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 403) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000011111111111100000000000000111111111111110000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001110011111000000000000000000111111111100000000000000000011111111110000000000000000011111111000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000001111111110000000000000000000011111111100000000000000000000011011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 404) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111100001110000000000000000111111000111000000000000000000001111111100000000000000000000011111100000000000000000000001111100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 405) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111100000000000000000111111111111000000000000000111111000011100000000000000011110000000110000000000000001110000000011000000000000000110000000000000000000000000011000000000000000000000000001100011000000000000000000000011111110000000000000000000001111111000000000000000000001111111100000000000000000001111111000000000000000000000111100000000000000000000000011100000100000000000000000001110000111000000000000000000111000111100000000000000000001111111110000000000000000000011111110000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 406) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001110000000111000000000000001111101110111100000000000000111111111111110000000000000001111111111111000000000000000010111100111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 407) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000001000000000000000001110000001111000000000000000111011111111100000000000000011111111111110000000000000001111111111110000000000000000011111100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 408) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111111100000000000000111111111111110000000000000111111000000000000000000000011111000000000000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000001100000001000000000000000000111001111110000000000000000001111111111000000000000000000011111110000000000000000000011111000000000000000000000011111000000000000000000000001110000000000000000000000000111000000000000000000000000001111111100000000000000000000111111110000000000000000000000111111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 409) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000001111111111111000000000000011111111111111110000000000011111111111111111000000000011111100000000000000000000011111000000000000000000000001110000000000000000000000000111000001110000000000000000011100111111100000000000000001111111111110000000000000000011111111110000000000000000011111111000000000000000000011111100000000000000000000001111000000000000000000000000111111110000000000000000000001111111100000000000000000000111111110000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 410) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000111111111100000000000000000111111111111000000000000000111110000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001100001110000000000000000000111111111100000000000000000001111111110000000000000000000111111110000000000000000000011111100000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000000111111110000000000000000000001111111000000000000000000000001111100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 411) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000011111111111100000000000000111111111111110000000000001111111111100011000000000000111111000000001100000000000111110000000000100000000000011110000000000000000000000001111000000000000000000000000011100111110000000000000000001111111111000000000000000000111111111100000000000000000011111111100000000000000000011111111100000000000000000001111100000000000000000000000111100000000000000000000000011110000100000000000000000000111111111000000000000000000011111111110000000000000000000111111110000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 412) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000011000000000000000000111110001110000000000000000011111111111000000000000000000110111111000000000000000000000000111100000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 413) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000001100000000000001110000000001110000000000000111000000001111000000000000011111011111111000000000000001111111111111100000000000000111111111111100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 414) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000011111111111000000000000000011111111100000000000000000011111000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000010000000000000000001110001111000000000000000000111111111100000000000000000001111111100000000000000000000111110000000000000000000000111100000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000001110000000000000000000000000111111111100000000000000000001111111110000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 415) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000001111111110000000000000000011111110000000000000000000011111000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000011000001000000000000000000000111111110000000000000000000011111110000000000000000000001111111000000000000000000001111100000000000000000000001111100000000000000000000001111000000000000000000000000111000000000000000000000000111110000100000000000000000011111111111000000000000000000111111111100000000000000000000000011100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 416) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000011111000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000001000000000000000000111000011100000000000000000011111111111000000000000000001111111111100000000000000000111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 417) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000111111111110000000000000001111111111000000000000000001111111000000000000000000011111100000000000000000000011111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110001100000000000000000000011111111000000000000000000000111111100000000000000000000111111100000000000000000000111111000000000000000000000011111000000000000000000000001111000000000000000000000000111111100000000000000000000001111111000000000000000000000000111110000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 418) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000001111111111000000000000000011111111111110000000000000111111000000111000000000000111100000000001000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000001100000000000000011100000011110000000000000000111111111111000000000000000001111111110000000000000000000011111100000000000000000000001111100000000000000000000001110000000000000000000000000111000000000000000000000000011100111111100000000000000001111111111100000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 419) begin
            pixels = 784'b0000000000000000000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000011000000000000000000000000001100000000000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000001000000000100000000000000001111000000010000000000000000111111000001000000000000000011101111101100000000000000000000001111110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 420) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011000011000000000000000000001100111100000000000000000000111111100000000000000000000011111100000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 421) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000010000000000000000000111000011100000000000000000011000001110000000000000000001100000110000000000000000001110000011000000000000000000111000011100000000000000000011101001110000000000000000001111111111000000000000000000111111111000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 422) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000011111111110000000000000000011111111011100000000000000111111100001110000000000000011100000000011000000000000011100000000001100000000000011100000000000000000000000001110000000000000000000000000110000000011000000000000000011100001111100000000000000000111111111110000000000000000011111111100000000000000000001111111100000000000000000000111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011110000001100000000000000000111111111110000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 423) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000011110000000000000000000000011111000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100111110000000000000000011111111111111110000000000001111111111111111000000000000000000000001111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 424) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000111111100000000000000000000111100100000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001111100000000000000000000000011111100000000000000000000000011111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000111100000000000000001111111111110000000000000000111111111111000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 425) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001111111000000000000000000000111111111110000000000000000011111111111000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 426) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111110000000000000000000111111111000000000000000000011111001100000000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000000110000000000000000000000000011100000000000000000000000000011000000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000110000111000000000000000000011111111100000000000000000000111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 427) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000001111100000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000001111110000000000000000000000111110000000000000000000000011100000000000000000000000111100000000000000000000000011110000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000001111100011111111000000000000111111111111111100000000000011111111111111110000000000000111111111111111000000000000001101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 428) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111110000000000000000011111111111000000000000000111111111111100000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111110000000000000000000000000111110000000000000000000000000111111000000000000000000000011111100000000000000000000001111110000000000000000000001110000000000000000000000001110000000000000000000000011110000000000000000000000011111000111100000000000000011111111111110000000000000000111111111111000000000000000011111111110000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 429) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000111001100000100000000000000011111111111111000000000000001111111111111100000000000000011111111111110000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 430) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011001100000000000000000000001111111111110000000000000000111111111111100000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 431) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001111111111111000000000000000111111111111110000000000000001111111111111000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 432) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011111000000000000000000000111111100000000000000000001111111110000000000000000001111100110000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011110000000000000000000000000111100000000000000000000000011110000000000000000000000000111000000000000000000000000111100000000000000000000000011000000000000000000000000111000000000000000000000000111000000000000000000000000011110111110000000000000000001111111111000000000000000000111111111100000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 433) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000001000000000000000111111111111111000000000000011111111111111100000000000001111111111111100000000000000111111111111100000000000000001101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 434) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000011111110000000000000000000011111000000000000000000000011110000000000000000000000011110000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011111100000000000000000000000111111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000001000000000000000000000000001100000000000000000000000001100000001100000000000000000111111111110000000000000000011111111110000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 435) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000011111100000000000000000000111111000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111110111100000000000000000001111111110000000000000000000001111110000000000000000000000111111000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000011110011110000000000000000000111111110000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 436) begin
            pixels = 784'b0000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000100000000000000000000000001111000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001111111111110000000000000000011111111111100000000000000000111010111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 437) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000011111111111000000000000000111111111111100000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000000111110000000000000000000000011111100000000000000000000000011111000000000000000000000000111000000000000000000000011110000000000000000000000011100000000000000000000000011110000000000000000000000011100000000000000000000000001110000000000000000000000001110000000011111000000000001111111111111111100000000000111111111111111100000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 438) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111111000000000000000001111111111110000000000000001111100000111000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000000111110000000000000000000000000111100000000000000000000000001111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000111000000000000000000000001100000000000000000000000011110000000000000000000000001111000000001111000000000000111111111111111110000000000001111111111111110000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 439) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111111111111000000000000000011111111111100000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 440) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000011111100000000000000000000011110110000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000000110000000000000000000000000111000000000000000000000000001111110000000000000000000000001111100000000000000000000001111000000000000000000000000111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000100000000000000000111000111111000000000000000011000111111100000000000000001111111111100000000000000000111111110000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 441) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111110000000000000000001111110011000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011110000000000000000000000000111100000000000000000000000011110000000000000000000000011100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000111100000000000000001111111111110000000000000000111111111110000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 442) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000001111111100000000000000000011111111110000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011110000000000000000000000000111111000000000000000000000001111110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001100001110000000000000000001111011111000000000000000000111111111000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 443) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111000011111110000000000000111111111111111000000000000011111111111111100000000000001111111110001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 444) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000100000000000000001111111111111111000000000000011111111111111100000000000000111100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 445) begin
            pixels = 784'b0000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000011000000000000011111111111111110000000000000111111111111111000000000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 446) begin
            pixels = 784'b0000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111100000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111000000000000000000000000111100000000000000000000000011110111111110000000000000011111111111111000000000000001111111111111100000000000000111111111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 447) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000001111110000000000000000000011111100000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000011110000000000000000000000000011000000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000011000011110000000000000000001111111111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 448) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111110000000000000000001111111111000000000000000001111100000100000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000011111000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011111100010000000000000000000111111111100000000000000000001111111110000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 449) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000011000000000000000110000000011100000000000000011000000001100000000000000001101111111110000000000000000111111111110000000000000000001100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 450) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000111111100000000000000000001111111111000000000000000001111000001110000000000000001110000000011000000000000000110000000000100000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001110000000000000000000000000011000000000000000000000000001110000100000000000000000000011111110000000000000000000000111110000000000000000000000011100000000000000000000000011100000000001000000000000001100000000011100000000000000111111111111100000000000000011111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 451) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000010000000000000000001100000001100000000000000000110000001110000000000000000010000111111000000000000000011111111111000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 452) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000001111111111111000000000000011111100000011100000000000011100000000000110000000000011100000000000001000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001110000000000000000000000000011000000110000000000000000001111001111000000000000000000011111110000000000000000000000111100000000000000000000000111000000000000000000000000011000000000000000000000000011100000001100000000000000000111111111110000000000000000011111111110000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 453) begin
            pixels = 784'b0000000000000000010000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000001100000000000000000000000001100000000000000000000000000100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000010000000000000011000000000011000000000000011000000000001100000000000001100000000000110000000000001110000000000011000000000000110001100000011000000000000011111111111111100000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 454) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000100000000000000001110000000110000000000000000110000000111000000000000000011000001111100000000000000001111111111110000000000000000011001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 455) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000011111111110000000000000001111111101111000000000000011111100000000100000000000011110000000000110000000000011110000000000110000000000011100000000000000000000000001100000000000000000000000000110000011000000000000000000011001111100000000000000000001111111100000000000000000000011111000000000000000000000011110000000000000000000000011100000000000000000000000011100000000011000000000000001110000111111100000000000000111111111111100000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 456) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111000000000000000000011111111111100000000000000111111100001111000000000000111100000000000110000000000011000000000000001000000000001100000000000000000000000000100000000000000000000000000011000000000000000000000000000110000000000000000000000000001111111100000000000000000000111111000000000000000000000111110000000000000000000011100000000000000000000000011110000000001100000000000000111111111111100000000000000001111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 457) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000011111111111100000000000000111111000000111000000000001111100000000000100000000001111000000000000000000000001111000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000000100000011000000000000000000011000111110000000000000000000111111100000000000000000000001111000000000000000000000001111100000000000000000000000111100000011111000000000000011000001111111100000000000000111111111111000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 458) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111111100000000000000011111111111111100000000000011111100000001110000000000011110000000000000100000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000000100000000000000000000000000011000000000000000000000000000011000000000000000000000000000111110000000000000000000000001111100000000000000000000001111000000000000000000000101111000000000000000000001111110000000000000000000001111100000001000000000000000111100000111110000000000000001111111111111000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 459) begin
            pixels = 784'b0000000000000000000000000000000000000000110000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000100000000000000001110000000010000000000000000110000000011000000000000000011000000001100000000000000011100000001110000000000000001110011111111000000000000000111111111111000000000000000011111100000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 460) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000001111111111100000000000000011111111111110000000000000011111100000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000110000000000000000000000000011100001100000000000000000000011111111000000000000000000001111111000000000000000000011111110000000000000000000111111100000000000000000000011110000000000000000000000001110000000000000000000000000110000000000000100000000000011110000011001111000000000000111111111111111000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 461) begin
            pixels = 784'b0000000000000000000000000000000000000000000000100000000000000000000000000011000000000000000000000000001000000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000010000000000000000111000000011000000000000000011000000001100000000000000001000000001110000000000000001111011111110000000000000000111111111111000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 462) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111111100000000000000001111000000110000000000000011110000000001100000000000001100000000000100000000000001100000000000010000000000000110000000000000000000000000001000000000000000000000000000110000000000000000000000000001100000110000000000000000000011111111000000000000000000000111111000011111100000000000111111111111111110000000000011111111111111000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 463) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011000000110000000000000000011000000010000000000000000001100000011000000000000000001100000001100000000000000000100011111100000000000000000011111111110000000000000000001111000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 464) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000111111110000000000000000011111111111100000000000000111111100000100000000000000111110000000000000000000000011000000000000000000000000001000000000000000000000000000110000000000000000000000000001100000000000000000000000000111110000000000000000000000011111000000000000000000011111100000000000000000000011111000000000000000000000011111111111110000000000000001111111111110000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 465) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000111111111111000000000000001111111111111110000000000001111111100011111100000000000111100000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000001110000000000000000000000000111111110000000000000000000001111111000000000000000000001111110000000000000000000011111110000000000000000000011111000000000000000000000001111000000000000000000000000111111111111111000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 466) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111111000000000000000011111111111110000000000000111111100000011000000000000111110000000000100000000000111100000000000010000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000001000000001100000000000000000011111111110000000000000000000011111110000000000000000000001111110000000110000000000001111100000001111100000000000111000111111111110000000000011111111111111100000000000001111111111100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 467) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111100000000000000001111111111111110000000000011111111111111111100000000011111111000000011110000000001111000000000000011000000001110000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000011111000000000000000000000000111111111100000000000000000000111111110000000000000000000011111100000000000000000000001110000000000000000000000001110000001110000000000000000111111111111000000000000000111111111111000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 468) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000100000000000000001111000000110000000000000001110000000011000000000000000110000000011100000000000000111000000001110000000000000011100000000110000000000000001111111110010000000000000000111111111111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 469) begin
            pixels = 784'b0000000000000000000000000000000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000100000000000000011100000000010000000000000001100000000011000000000000000110000000011100000000000000000000000011110000000000000000000000001110000000000000001011111111110000000000000000111111111110000000000000000001000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 470) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011101000110000000000000000001100000010000000000000000001110000011000000000000000000110000011000000000000000000010000001100000000000000000011000001100000000000000000011001111000000000000000000001111101100000000000000000001111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 471) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111100000000000000000000111111110000000000000000000111100011100000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111110000000000000000000000011111000000000000000000000001111100000000000000000000000111100000000000000000000000011100001000000000000000000011100001110000000000000000001110000111000000000000000000111001111100000000000000000011111111100000000000000000001111111110000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 472) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000011000000000000000000011100001110000000000000000000111111111000000000000000000011111111100000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 473) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000001111110000000000000000000011111111100000000000000000011111111110000000000000000011111000011000000000000000001111000001100000000000000000111000000000000000000000000011100000000000000000000000001110001100000000000000000000111111110000000000000000000011111111000000000000000000000111111100000000000000000000111111100000000000000000000011100000000000000000000000011110000000000000000000000000111000110000000000000000000011111111000000000000000000000111111100000000000000000000001111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 474) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000110000000000000000011100000111000000000000000011110000011100000000000000001110001111110000000000000000111111111111000000000000000001111111111100000000000000000111111111110000000000000000000111000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 475) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011111000000000000000000000011111111000000000000000000011111111100000000000000000011110011110000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000001110111000000000000000000000111111110000000000000000000001111111000000000000000000000111111000000000000000000000111100000000000000000000000011100000000000000000000000001110000011000000000000000000111101111100000000000000000001111111110000000000000000000111111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 476) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000111000000000000000011100000011100000000000000001110000001110000000000000000111111111110000000000000000001111111111000000000000000000111111111100000000000000000001110000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 477) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000110000000000000000011000000111000000000000000011100000011100000000000000001110000111110000000000000000111111111110000000000000000011111111111000000000000000001111111111000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 478) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000011000000000000000000111000011100000000000000000011111111110000000000000000001111111110000000000000000000111111111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 479) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000111111111000000000000000000111111111100000000000000000011111111110000000000000000011100000110000000000000000011100000000000000000000000001110000000000000000000000000111000010000000000000000000011111111100000000000000000001111111110000000000000000000011111110000000000000000000001111100000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000100000000000000000111000011110000000000000000011111111111000000000000000001111111111000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 480) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111100000000000000000011111111110000000000000000011111111111000000000000000001111000000000000000000000000111000000000000000000000000111110000000000000000000000001111000011000000000000000000111111111100000000000000000001111111111000000000000000000111111111000000000000000000001111111000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001110000011110000000000000000111100011111000000000000000011111111111100000000000000001111111111000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 481) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111110000010000000000000000011110000011100000000000000001111000011110000000000000001111000001111000000000000000111100001111100000000000000011110000111110000000000000011111111111111000000000000001111111111111000000000000000111111111111100000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 482) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000111111111111000000000000000111111111111100000000000001111111100001110000000000001111110000000011000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000000011111110000000000000000000000111111000000000000000000000011111100000000000000000000011111110000000000000000000011111000000000000000000000001111000000000000000000000000111000000000000000000000000011100001111000000000000000001111011111100000000000000000011111111110000000000000000000111111110000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 483) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111000000000000000000111111111110000000000000000111111111111000000000000001111111111111100000000000000111111000001110000000000000011110000000010000000000000001111000000000000000000000000111000000000000000000000000001110011110000000000000000000111111111100000000000000000011111111110000000000000000011111111111000000000000000011111110000000000000000000001111100000000000000000000000111110000111000000000000000001111111111100000000000000000111111111110000000000000000000111111111100000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 484) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000111111000000000000000000000111111110000000000000000001111111111100000000000000000111111111110000000000000000111111000110000000000000000011111000000000000000000000001111000000000000000000000000111111000000000000000000000001111110000000000000000000000111111000000000000000000000111111100000000000000000000111111100011000000000000000011111000011100000000000000001111000011110000000000000000111111111111000000000000000001111111111100000000000000000111111111100000000000000000001111111100000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 485) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000001100000000000000000011110011111000000000000000001111111111100000000000000000111111111100000000000000000000111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 486) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000011111100000000000000000000011111111000000000000000000011110011000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111101100000000000000000000011111111000000000000000000000111111000000000000000000000001111100000000000000000000000111000000000000000000000000111000000000000000000000000011000000110000000000000000001110000111000000000000000000111000111000000000000000000001111111000000000000000000000011111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 487) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000011100000000000000011100000011110000000000000011110000001111000000000000001111001111111000000000000000111111111111100000000000000011111111111110000000000000000111000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 488) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000010000000000000000011110000011100000000000000001111000001110000000000000000111100001111000000000000000001111111111000000000000000000111111111100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 489) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001110000000111000000000000000111111110111100000000000000011111111111100000000000000000111111111110000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 490) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111110000000000000000000111111111000000000000000000111111111100000000000000000111111000000000000000000000011111000000000000000000000001111000000000000000000000000111001110000000000000000000011111111000000000000000000001111111110000000000000000000011111111000000000000000000011111111000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000011100000000000000011110001111110000000000000000111111111111000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 491) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000011111111000000000000000000011111111100000000000000000011111100010000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100011100000000000000000000111111110000000000000000000011111110000000000000000000001111110000000000000000000000111100000000000000000000000111100000000000000000000000111100001110000000000000000011100011111000000000000000001111111111100000000000000000011111111100000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 492) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011110000001000000000000000001111000001100000000000000000111000001111000000000000000111111111111000000000000000001111111111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 493) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000001100000000000000001110000001110000000000000000111000001111000000000000000001111111111100000000000000000011111111100000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 494) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000100000000000000000011100000111000000000000000011110000111100000000000000001111000011110000000000000000111111111110000000000000000011111111110000000000000000000111111111000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 495) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000011111111000000000000000000011111111110000000000000000011111111111000000000000000011111000001100000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011111111000000000000000000000111111100000000000000000000011111100000000000000000000001111110000000000000000000001111100000000000000000000001111000011000000000000000000111001111100000000000000000111111111110000000000000000001111111111000000000000000000111111110000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 496) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111111000000000000000000011111111110000000000000000011111111111000000000000000011110000001100000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000000111100000000000000000000000011111110000000000000000000000111111000000000000000000000111111100000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000011100001000000000000000000001111111110000000000000000000011111110000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 497) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000011111111111100000000000000011111000011111000000000000111110000000001100000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000001100000001000000000000000000110000111100000000000000000011111111110000000000000000000111111111000000000000000000000111111000000000000000000000000111000000000000000000000000011111110000000000000000000001111111000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 498) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111110000000000000000001111100011100000000000000001110000000100000000000000001110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000011100000000000000000110000111110000000000000000011111111100000000000000000000111110000000000000000000000001110000000000000000000000001100000000000000000000000000110000000001110000000000000011100111111110000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 499) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000001111000000000000000110000111111110000000000000011111111111111000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 500) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110001111000000000000000000001111111000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 501) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000111111110000000000000000001111100001000000000000000001111000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000001000000000000000011100000011100000000000000001110001111100000000000000000111011111100000000000000000001111111100000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000000111111111100000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 502) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000011110000000000000000000000001110000000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001111111110000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 503) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111000000000000000011111110001100000000000000011110000000010000000000000011110000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000001110001100000000000000000000111111110000000000000000000001111110000000000000000000000111100000000000000000000000011100000000000000000000000111100000011110000000000000111100000111110000000000000011111111111110000000000000011111111111100000000000000001111111110000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 504) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000001111111110000000000000000001111100001000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001100011110000000000000000000111111110000000000000000000011111110000000000000000000000111100000000000000000000000111100000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000111111000000000000000011111111111100000000000000001111111111000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 505) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000001000000000000001111000000011110000000000000011111111111100000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 506) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000111111010000000000000011111111110000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 507) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111000000000000000000111100000010000000000000000111100000001000000000000000111000000000100000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000001100000000000000000000000000110000011100000000000000000011111111000000000000000000000111111000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000011000000110000000000000000011111111111000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 508) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000001111100000000000000001110111111110000000000000000011111110000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 509) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000001111110000000000000011111111111111100000000000001111111000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 510) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000111111111000000000000000001111110001110000000000000001111000000011000000000000011110000000011100000000000001110000000001100000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000010000000000000000000111111111100000000000000000001111111100000000000000000000011110000000000000000000000111100000000000000000000000111000000000000000000000000111000000000000000000000000111000000000111000000000000001111111111111110000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 511) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000111111000000000000000000000111111110000000000000000000111110011100000000000000000111100000110000000000000000011100000011000000000000000011100000001100000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000010000000000000000000001110111100000000000000000000111111100000000000000000000001111100000000000000000000000111100000000000000000000000011100000000000000000000000011111111100000000000000000001111111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 512) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001110000000011100000000000000111000011111110000000000000001111111111110000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 513) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000011111111000000000000000000011110000110000000000000000011110000001000000000000000001110000001100000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000110000000000000000000111001111000000000000000000001111111000000000000000000000111110000000000000000000000011110000000000000000000000001110000000000000000000000001110011100000000000000000000110011110000000000000000000011111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 514) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111110000000000000000011110000011000000000000000011110000001100000000000000011100000001100000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011000000000000000000000000011100001111000000000000000001100111111100000000000000001100111111100000000000000000111111110000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 515) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000111110000000000000000000000111100000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000001111111110111000000000000000011111110000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 516) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000111100000000000000001110011111110000000000000000111111111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 517) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111111000000000000000001111000001100000000000000001111000000110000000000000001110000000011000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110001110000000000000000000011111111000000000000000000000111111000000000000000000000011110000000000000000000000011110000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110011111110000000000000000011111111110000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 518) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000001111100000000000000000000001111000000000000000000000001111100000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000000111000000011110000000000000011111111111111000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 519) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111111000000000000000111111111111110000000000000011110000001110000000000000011100000000010000000000000011100000000000000000000000001100000000000000000000000001110000001110000000000000000111000011111000000000000000011111111111100000000000000000111111111000000000000000000001111110000000000000000000000111100000000000000000000000111100000000000000000000000111100011000000000000000000011100111100000000000000000011111111110000000000000000000111111110000000000000000000001111110000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 520) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000001110000000000000111000000011111000000000000011100000111111000000000000001100111111110000000000000001111111111110000000000000001111111000010000000000000000111100000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 521) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000111111110000000000000000001111111111100000000000000001111110001111100000000000000111000000011110000000000000111000000000111000000000000111000000000000000000000000011100000100000000000000000011100011111000000000000000001111111111000000000000000000011111110000000000000000000001111110000000000000000000000111100000000000000000000000111100010000000000000000001111100111100000000000000000111111111110000000000000000111111111110000000000000000001111111110000000000000000000000011110000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 522) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001111000001110000000000000001111000111111100000000000001111111111111100000000000001111111111111000000000000001111111100000000000000000000111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 523) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000001111111111100000000000000001111111111110000000000000001111000000111100000000000001110000000011100000000000001110000000000010000000000000111000000000000000000000000111000000000000000000000000011000001110000000000000000001111111111100000000000000000111111111100000000000000000011111110000000000000000000000111100011000000000000000000111100111110000000000000000111111111110000000000000000011111111110000000000000000001111111100000000000000000000111111100000000000000000000001111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 524) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000110000000000000000111100000111000000000000000111000000111100000000000000011101111111110000000000000011111111111110000000000000001111111111110000000000000000111100011110000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 525) begin
            pixels = 784'b0000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000100000000000000000001110000111000000000000000000110000111000000000000000000111011111000000000000000000011111111000000000000000000011111111000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 526) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000001111111111110000000000000011111000001111100000000000001110000000001111000000000001110000000000011000000000001111000000000000000000000000110000001110000000000000000011000011111000000000000000001100111111000000000000000000111111110000000000000000000001111100000000000000000000001111000000000000000000000001111000000000000000000000001111000011000000000000000000111000111110000000000000000011111111111000000000000000000111111100000000000000000000000111100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 527) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000010000000000000000011110000111100000000000000001110001111110000000000000001111111111110000000000000000111111111110000000000000000011111000010000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 528) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111111100000000000000000011111111111000000000000000011111111111110000000000000011110000000111000000000000001110000000011100000000000000110000000000110000000000000011000000000000000000000000011100000110000000000000000001110001111000000000000000000011101111000000000000000000001111111000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001111011100000000000000000001111111110000000000000000000111111111000000000000000000011111111000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 529) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111110000000000000000011111101111100000000000000011110000001111000000000000011110000000011100000000000001110000000000110000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000110000000000000000000011111111000000000000000000001111111100000000000000000000011111000000000000000000000001111000000000000000000000001110000000000000000000000000111001110000000000000000000011111111000000000000000000001111111000000000000000000000011111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 530) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000010000000000000001111000000111100000000000001111000000111110000000000001111000001111110000000000001111111111111110000000000000111111111111110000000000000111111111111110000000000000111111100001110000000000000011111000000011000000000000001110000000001100000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 531) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001111111111000000000000000011111111111111000000000000011111000001111110000000000011110000000000111000000000011110000000000001000000000001110000011000000000000000001110000111100000000000000000111001111110000000000000000011111111100000000000000000001111111000000000000000000000011111000000000000000000000001110000100000000000000000001110000111000000000000000001110001111000000000000000000111111111000000000000000000011111111000000000000000000000111111000000000000000000000001111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 532) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001100001110000000000000000001111111111000000000000000000111111111000000000000000000111110011000000000000000000011100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 533) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000111000000000000000001110000011100000000000000000111000111110000000000000000111101111110000000000000000011111111110000000000000000001111111110000000000000000000111111000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 534) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000001111111100000000000000000001111111111000000000000000011111000011100000000000000011110000001110000000000000011100000000011000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000011100000000000000000001100111110000000000000000000111111110000000000000000000001111100000000000000000000000011100000000000000000000000011100000100000000000000000011100001111000000000000000001110001111100000000000000000111111111000000000000000000011111111000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 535) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000111111111000000000000000000111100011110000000000000000111000000111100000000000000111000000001100000000000000011000000000000000000000000001100000011000000000000000000111000111100000000000000000011101111100000000000000000000111111000000000000000000000001111000000000000000000000000111000000000000000000000000111000110000000000000000000111000111000000000000000000111001111100000000000000000011111111100000000000000000001111111000000000000000000000011111000000000000000000000000011000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 536) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000010000000000000011000000000111000000000000011100000001111100000000000001111001111111100000000000001111111111111100000000000000111111111111100000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 537) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110011111100000000000000000111111111110000000000000000111111110011000000000000000011111100000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 538) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000110000000000000000000111011111100000000000000000011111111000000000000000000011111100000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 539) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000001111111100000000000000000001111000110000000000000000000110000011000000000000000000110000000000000000000000000011000000000000000000000000000110000000000000000000000000011100000000000000000000000000111100000000000000000000000001111100000000000000000000000001111111111000000000000000000001111111000000000000000000000011111000000000000000000000011110000000000000000000000011110000000000000000000000011100000000000000000000000001111100000000000000000000000111111111101000000000000000000001111111110000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 540) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000111000000000011111111111111111111000000000111111111111011111100000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 541) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000011111100000000000000000000011110110000000000000000000011100010000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000000111000000000000000000000000011111000000000000000000000000011111110000000000000000000000011111110000000000000000000000011111000000000000000000000011111000000000000000000000111110000000000000000000001111100000000000000000000001111000000100000000000000000111100000111000000000000000011111111111000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 542) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000111111000000000000000000001111110000000000000000000001111000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000011110000000000000000000000000011111000000000000000000000000111111000000000000000000000000111111100000000000000000000000011110000000000000000000000111111000000000000000000001111100000000000000000000001111000000000000000000000000111000000000000000000000000011111000000000000000000000000011111111110000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 543) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000111000000000000000000000000011111111111110000000000000000001111111111100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 544) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111100000000000000000111110000010000000000000000111100000000000000000000000111100000000000000000000000011000000000000000000000000011100000000000000000000000000110000000000000000000000000001100000000000000000000000000111100000000000000000000000001111100000000000000000000000001111111111000000000000000000000111111100000000000000000000001111100000000000000000000011110000000000000000000000111100000000000000000000000111000000000000000000000000011100000000000000000000000001111111111110000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 545) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000111111100000000000000000000111111100000000000000000000111100000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001111100000000000000000000000011111111110000000000000000000011111111000000000000000000000001111000000000000000000000111110000000000000000000001111100000000000000000000001111000000000000000000000000111000000000000000000000000011111111110000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 546) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111111111111111110000000000011111111111111111110000000000000000111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 547) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001111000000000000000000000000111111111110000000000000000000111111111111000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 548) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111111100000000000000000000000111111111100000000000000000000001111111100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 549) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011111111111100000000000000001111111111110000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 550) begin
            pixels = 784'b0000000000000000000000000000000000000000000100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000011000011110000000000000000001111111111111000000000000000001110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 551) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000001111111000000000000000000000111111100000000000000000000111000110000000000000000000111100001000000000000000000011100001000000000000000000001111000100000000000000000000111100000000000000000000000001111110000000000000000000000011111111111000000000000000000111111111110000000000000000000011111110000000000000000000000011110000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111101011000000000000000000011111111110000000000000000000111111110000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 552) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000111111111000000000000000000111000000000000000000000000111000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000001110000011000000000000000000011111111100000000000000000000011111100000000000000000000000111000000000000000000000000110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000110000000000000000000111111110000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 553) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000111110000000000000000000000111000100000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000001111110000000000000000000000011111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000110000000000000000000011111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 554) begin
            pixels = 784'b0000000000000000000000000000000000000000001000000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000000111111111111100000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 555) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000011111100000000000000000000001100010000000000000000000001100001000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000000110000000000000000000000000011100000000000000000000000000111110010000000000000000000000111111000000000000000000000000111000000000000000000000000111000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000000011000011000000000000000000001111111000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 556) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000111110000000000000000000000111101100000000000000000000011100110000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000000110000000000000000000000000011100000000000000000000000000111000000000000000000000000001111100000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011111110000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 557) begin
            pixels = 784'b0000000000011000000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000011100000000000011110000111111110000000000000111111111111110000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 558) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000000111100000000000000000000000001111111000000000000000000000000111111110000000000000000000000001111111000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 559) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000000111000000000000000000000000001111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 560) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000011111111100000000000000000011100000010000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000001111000000000000000000000000001111000000000000000000000000011111110000000000000000000000001111000000000000000000000001110000000000000000000000011100000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011110000011000000000000000000111111111110000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 561) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000011111111100000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000001000000000000000000000000000110000000000000000000000000001100000000000000000000000000011100000000000000000000000000111111110000000000000000000000111110000000000000000000000011100000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000000111100000000000000000000000001111111100000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 562) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000111111111110000000000000000111111111111100000000000000111111111111111000000000000111111110001111100000000000011111000000111100000000000011111000000001100000000000001111000000000000000000000001111111100000000000000000000111111111000000000000000000001111111100000000000000000000111111100000000000000000000001111100000000000000000000000111100011100000000000000000011110111110000000000000000001111111111000000000000000000111111111100000000000000000011111111100000000000000000001111111000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 563) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000001111100000001000000000000000111110000001110000000000000111111110001111100000000000011111111111111110000000000011111111111111110000000000001111111111111110000000000000111111111111100000000000000011110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 564) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000001111111110000000000000000011111111111000000000000000111111111111100000000000000111111111101100000000000000111111100000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000000111111110000000000000000000001111111100000000000000000000111111110000000000000000000011111110000000000000000000001111110000000000000000000001111110000000000000000000000111110000000000000000000000011111111110000000000000000001111111111111000000000000000111111111111100000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 565) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011111000000000000000000000011111100000000000000000000001111100000000000000000000001111100000000000000000000001111110000000000000000000000111110000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000011110000000000001111100111111111000000000000011111111111111100000000000001111111111111100000000000000111111111110000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 566) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000111111111110000000000000000111111111111100000000000001111111110111100000000000001111110000011100000000000001111100000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000011111111000000000000000000001111111110000000000000000000011111111000000000000000000001111111000000000000000000000111110000000000000000000000111100000000000000000000000011110000000000000000000000011111000111000000000000000000111111111110000000000000000011111111111000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 567) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000001111100000001000000000000000111100000001110000000000000111110000011111000000000000011110000011111000000000000001111100011111000000000000000111111111111000000000000000011111111110000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 568) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000100001111000000000000000000010001111000000000000000000001000111100000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000010000000000000000001110000011100000000000000001111000011110000000000000000111111001110000000000000000011111111111000000000000000001111111111000000000000000000111111111100000000000000000011000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 569) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000011000000000000000111110000011100000000000000011110000011110000000000000001111111111111000000000000001111111111111000000000000000111111111111100000000000000011111111111100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 570) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000111111110000000000000000001111111111000000000000000011111111111000000000000000111111100001000000000000000111111100000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000001111100000000000000000000000111110011110000000000000000011111111110000000000000000001111111111000000000000000000011111111000000000000000000000011111000000000000000000000001111000000000000000000000000111100111100000000000000000011111111110000000000000000001111111110000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 571) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000011100000000000001110000000001110000000000001111000000001111000000000000111100000000111100000000000111110000000111100000000000011111111110011100000000000001111111111111110000000000000111000001111110000000000000010000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 572) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111110000000000000000001111111111000000000000000001111111111110000000000000011111110000010000000000000001111100000000000000000000001111000000000000000000000000111000000000000000000000000111100111000000000000000000011111111110000000000000000001111111110000000000000000000011111110000000000000000000001111110000000000000000000000011110000000000000000000000011110000100000000000000000001111000111000000000000000000111111111110000000000000000011111111110000000000000000000111111110000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 573) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000111110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000001111100000000000000000000000111110000011100000000000000111110000011110000000000000011110000001111000000000000011111110011111000000000000001111111111111000000000000000111111111111000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 574) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000111111111111100000000000000011111111111110000000000000011111111111111000000000000011111111111111000000000000011111000011110000000000000001110000000000000000000000001111000000000000000000000000111000000100000000000000000111100111110000000000000000011111111111000000000000000000111111111100000000000000000011111111000000000000000000000111110000000000000000000000111110000000000000000000000011100000100000000000000000011111111111000000000000000011111111111100000000000000000111111111100000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 575) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000011111111111100000000000000111111111111111000000000000111111111111111100000000000111110111111111100000000000111110001111111100000000000011100000000110000000000000011100000000000000000000000001100000000000000000000000000110000000110000000000000000011100111111100000000000000001111111111110000000000000000011111111100000000000000000000111111100000000000000000000000111000000000000000000000000011100000000000000000000000001110000011000000000000000000111111111111000000000000000001111111111100000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 576) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000001000000000000000111100000001110000000000000011110000011111000000000000001111100011111100000000000000111111111111110000000000000011111111111110000000000000001111111111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 577) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000011111111100000000000000000111111111110000000000000000111111111111100000000000000111111101111100000000000000111111000011100000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011111000000000000000000000000111111000000000000000000000001111110000000000000000000001111111000000000000000000000111111000000000000000000000111110000000000000000000000001110000000000000000000000000111111111000000000000000000011111111110000000000000000000011111111000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 578) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000001111111111110000000000000001111111111111000000000000011111111111111110000000000011111111111111110000000000011111011111111100000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011111111110000000000000000000111111111000000000000000000011111111000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000000011111000010000000000000000001111111111100000000000000000001111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 579) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011111000000000000000000000111111000000000000000000000111111100000000000000000000011111100000000000000000000011111110000000000000000000001111110000000000000000000001111110000000000000000000000111110000000000000000000000111111000000000000000000000011111100000000000000000000001111100000000000000000000001111110000000000000000000000111110000000000000000000000011111000001111110000000000001111111111111111000000000000111111111111111100000000000011111111111111100000000000001111111110000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 580) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000011111111111000000000000000111111111111110000000000000111111111111110000000000000011111111111100000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000000111100100000000000000000000011111111000000000000000000001111111100000000000000000000011111100000000000000000000001111100000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001111001111000000000000000000111111111110000000000000000001111111110000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 581) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111110000000000000000011111111111100000000000000011111111111110000000000000111111111111110000000000000011110000001110000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001111111110000000000000000000111111111000000000000000000001111111000000000000000000000111111000000000000000000000111110000000000000000000000001111000000000000000000000000111111100110000000000000000001111111111000000000000000000011111111100000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 582) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111111100000000000000111111111111111000000000000111111111111111100000000000111111111111111111000000000011111111000000111100000000001111110000000000100000000000111111000000000000000000000011111111110000000000000000000111111111100000000000000000001111111111000000000000000000111111111100000000000000000011111111111000000000000000001111111111110000000000000000111111111111000000000000000011111111111100000000000000000111111111111000000000000000001111111111000000000000000000001111111000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 583) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111000000000000000000000011111100000000000000000000011111100000000000000000000001111110000000000000000000001111110000000000000000000000111111000001100000000000000111111000001111000000000000111111100000111100000000000011111100000111110000000000011111110000111111000000000001111111111111111100000000000111111111111111100000000000011111111111111110000000000000111111111111110000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 584) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000111111111111100000000000001111111111111111100000000001111111110000011110000000000111110000000000010000000000001111110000000000000000000001111111110000000000000000001111111111100000000000000001111111111100000000000000000111111000000000000000000000011111111000000000000000000000111111100000000000000000000001111110000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 585) begin
            pixels = 784'b0000000000000000000000000000000000000000000111100000000000000000000000111110000000000000000000000011111000000000000000000000011111100000000000000000000011111100000000000000000000001111110000000000000000000001111110000000000000000000001111110000000000000000000000111110000000000000000000000111111000000000000000000000011111000000000000000000000011111100000000000000000000011111100000010000000000000001111100000011110000000000001111110000011111100000000000111111111111111110000000000111111111111111110000000000011111111111111110000000000000111111111111110000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 586) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010000000000000001111111111111110000000000001111111111111111110000000000111111111111111111000000000011110000000000011100000000000111111110000000010000000000011111111100000000000000000111111111110000000000000000011111111111000000000000000011111100000000000000000000001111100000000000000000000000111100011111000000000000000001111111111110000000000000000011111111111000000000000000000111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 587) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000001111110000000000000000000001111111000000000000000000000111111000000000000000000000111111000000000000000000000111111000000000000000000000011111100000000000000000000011111100000000000000000000001111110000000000000000000001111110000011110000000000001111110000111111100000000000111111001111111110000000000111111111111111110000000000011111111111111110000000000001111111111111100000000000000111111111000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 588) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000001111100000000000000000000000111110000000000000000000000111111000000000000000000000011111000000000000000000000001111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000001111100000111000000000000000111110000111110000000000000011111000111111000000000000011111000011111000000000000001111111111111100000000000001111111111111100000000000000111111111111100000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 589) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000001111111111110000000000000001111111111111100000000000001111110000111111000000000001111100000001111100000000000111100000000001100000000000011111011100000000000000000001111111110000000000000000000011111111100000000000000000011111111100000000000000000011111110000000000000000000011111001000000000000000000011111111110000000000000000000111111111100000000000000000011111111100000000000000000000011111100000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 590) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000110000000000000000011110000111100000000000000011111000111110000000000000001111000011110000000000000001111111111111000000000000000111111111111000000000000000111111111110000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 591) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000011111111110000000000000000111111111111100000000000000111111111111110000000000000111111110011111100000000000011111100000111110000000000011111000000001111000000000001111100000000011100000000000011111111110000000000000000001111111111000000000000000000011111111100000000000000000011111111110000000000000000001111111111000000000000000001111111100000000000000000000111110111000000000000000000011111111100000000000000000001111111111000000000000000000011111111100000000000000000000111111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 592) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000111110000000000000000000000111111000000000000000000000111111100000000000000000000111111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111110000000000000000000001111110000000000000000000001111110000000000000000000001111111001111000000000000001111111001111100000000000000111111001111110000000000000111111001111111000000000000011111111111111100000000000001111111111111100000000000000011111111111100000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 593) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000011111000000000000000000000011111110000000000000000000001111110000000000000000000001111110000000000000000000001111111000000000000000000001111111000000000000000000000111111000000000000000000000111111100000000000000000000011111100000000000000000000011111100000000000000000000001111100000000000000000000001111110000011000000000000000111110000111110000000000000111111000111111000000000000111111100111111100000000000011111111111111100000000000001111111111111100000000000000011111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 594) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111111111000000000000000111111111111111000000000000011111111111111110000000000001111111111111111100000000000111110000000111111000000000011111000000000111110000000000111111111000001110000000000011111111110000010000000000011111111111000000000000000001111111111000000000000000001111111110000000000000000000111110000111000000000000000001111111111110000000000000000111111111111000000000000000001111111111100000000000000000011111111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 595) begin
            pixels = 784'b0000000000000000000000000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111100000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000001111100000000000000000000001111100000110000000000000000111110000111100000000000000111110000111110000000000000111110000111111000000000000111111100111111000000000000011111111111111000000000000000111111111111000000000000000001000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 596) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000111100000000000000000000000111110000000000000000000000111111000000000000000000000011111000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000001111100000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000011111000111000000000000000011111000011110000000000000011111111111111000000000000011111111111111000000000000001111111111111100000000000000111111111111100000000000000011111111101000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 597) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111000000000000000000000111111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000001111100000000000000000000001111110000000000000000000001111110001110000000000000001111111001111000000000000000111111001111100000000000000111111101111110000000000000111111111111111000000000000111111111111111000000000000011111111111111000000000000000111111111111000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 598) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111100000000000000000000001111110000000000000000000001111110000000000000000000000111111000000000000000000000111111000000000000000000000111111000000000000000000000111111000000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000001111100000110000000000000001111110000111100000000000000111110000111110000000000000111111011111111000000000000111111111111111000000000000011111111111111000000000000001111111111111000000000000000011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 599) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000011111000000000000000000000011111001110000000000000000011111000111100000000000000001111000111100000000000000001111111111110000000000000001111111111100000000000000000011111111100000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 600) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001111111111111100000000000001111111111111111000000000001111111111111111110000000000111111000000001111100000000011110000000000001100000000000111000000000000000000000000001110000000000000000000000000111111111100000000000000000001111111111000000000000000000111111111100000000000000001111111111100000000000000000111111110000000000000000000111111000000000000000000000011111111000000000000000000001111111111000000000000000000011111111100000000000000000001111111110000000000000000000011111110000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 601) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111111000000000000000000011111111100000000000000000001111111111000000000000000001111000111000000000000000000111000000100000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000011111111110000000000000000000111111111000000000000000000001111111000000000000000000000111111000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000000011110001100000000000000000001111111111000000000000000000111111111000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 602) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000111110000000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111111111000000000000000000011111111111100000000000000000111111111111000000000000000000111111111100000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 603) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000111111100000000000000000000011111111100000000000000000001111111111011110000000000000110000111111111000000000000011000000111111000000000000000110000001111000000000000000011100000000000000000000000000111011100000000000000000000011111111000000000000000000001111111100000000000000000001111111110000000000000000000111111110000000000000000000111110000000000000000000000011110000000000000000000000001110000000000000000000000000011100001110000000000000000001111111111100000000000000000011111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 604) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011110000000000000000000000001111000000000000000000000001111100000000000000000000001111100000000000000000000001111110000000000000000000001111110000000000000000000001111110000000000000000000000111111000000000000000000000111111000000000000000000000111111000000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000000011110000000000000000000000001111111001100000000000000000011111111111111000000000000000111111111111100000000000000001111111111110000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 605) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111111100000000000000011111111111111000000000000011111100001111100000000000011110000000011110000000000001110000000000010000000000000111000000000000000000000000111100000000000000000000000011110000000111000000000000000111111011111100000000000000001111111111110000000000000000011111111110000000000000000000011111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111111101111000000000000000001111111111100000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 606) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000001111110000000000000000000000011111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000011110000000000000000000000001111111111111100000000000000111111111111110000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 607) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000001111000000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111110000000000000000000000111110000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000000111100011111110000000000000011111111111111100000000000000111111111111100000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 608) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000001111111111111100000000000001111111111111110000000000001111110001111110000000000001111100000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001111111111110000000000000000011111111111100000000000000000111111111100000000000000000001111111000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111100001111000000000000000011111111111110000000000000000111111111111000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 609) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111110000000000000000000111111111000000000000000000011111111000000000000000000001111111000000000000000000001111111100000000000000000001111111100000000000000000001111111000000000000000000001111111000000000000000000001111111000000000000000000001111111000000000000000000001111111000000000000000000000111111000000000000000000000011111000000000000000000000001111000000000000000000000000111110000000000000000000000011111111111111111100000000000111111111111111110000000000001111111111111111000000000000000101110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 610) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111111110000000000000001111111111111100000000000001111111111111110000000000001111111111111111000000000000111111000000000000000000000011110000000000000000000000011111000000000000000000000000111110000000000000000000000011111111111000000000000000000111111111100000000000000000000111111110000000000000000000011111100000000000000000000011111100000000000000000000001111000000000000000000001100111100000000000000000000011111111111111100000000000000011111111111110000000000000000011111111111000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 611) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000111111111111100000000000000111111111111111000000000000011111100111111100000000000011111000000001100000000000001111000000000000000000000000111100000000000000000000000001111000000000000000000000000111110000000000000000000000001111110000000000000000000000011111111000000000000000000000011111110000000000000000000001111111000000000000000000000111111100000000000000000000111111100000000000000000000111111011100000000000000000011111111111000000000000000000111111111110000000000000000011111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 612) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000011111100000000000000000000011111110000000000000000000001111111000000000000000000000111111000000000000000000000111111000000000000000000000011111000000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000000111110000110000000000000000011110001111111000000000000001111111111111100000000000000111111111111110000000000000001111111111110000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 613) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111000000000000000011111111111110000000000000011111110111111100000000000011111000000011110000000000011110000000000010000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000001111100001100000000000000000001111111111000000000000000000011111111100000000000000000011111111000000000000000000001111100000000000000000000001111000000000000000000000000111111111111110000000000000001111111111111000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 614) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111000000000000000001111111111111000000000000000111000000011100000000000000111100000000111000000000000011100000000000000000000000000110000000000000000000000000111000000000000000000000000011110000000000000000000000000111111111000000000000000000001111111100000000000000000000011111110000000000000000000011111100000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000110000000000000000001111111111100000000000000000011111111110000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 615) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000011111000000000000000000000011111100000000000000000000011111100000000000000000000111111100000000000000000000011111100000000000000000000011111100000000000000000000111111100000000000000000000011111100000000000000000000011111000000000000000000000011111000000000000000000000011111000000000000000000000001111111111111111110000000000011111111111111111000000000000111111111111111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 616) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111111111000000000000000000011111111110000000000000000001111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 617) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000011111000000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000001111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011110001111111110000000000001111111111111111000000000000011111111111111000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 618) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000001111111110000000000000000011111111111100000000000000001111110011111000000000000001111000111111100000000000000111000011111111000000000000011000000011111100000000000001100000000011110000000000000111000000000111000000000000011111111110000000000000000000111111111100000000000000000011111111100000000000000000001111111100000000000000000001111111000000000000000000000111110000000000000000000000011110000000100000000000000001111111011111100000000000000011111111111110000000000000000111111111111000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 619) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000001111111110000000000000000001111111111100000000000000001111000111111000000000000000111000001111100000000000000111000000111110000000000000011100000000011000000000000001110000000000000000000000000111000000000000000000000000001100000110000000000000000000111111111100000000000000000001111111110000000000000000000011111110000000000000000000001111100000000000000000000000111000000000000000000000000011100000000000000000000000001111110000000000000000000000111111111000000000000000000001111111110000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 620) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000111111111111111000000000000111111111111111110000000000011111111111111111000000000011111100001111111100000000001111000000000111110000000001111100000000000000000000000111110000000000000000000000001111111111100000000000000000111111111110000000000000000001111111111000000000000000000001111111100000000000000000000111111000000000000000000000111110000000000000000000000111110000000000000000000000011111000001100000000000000001111101111111000000000000000011111111111100000000000000000111111111100000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 621) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111000000000000000000000111111100000000000000000000111111100000000000000000001111111100000000000000000001111111000000000000000000001111111000000000000000000000111111000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000000111110000000000000000000000001111111111110000000000000000011111111111110000000000000000111111111111000000000000000000111111111100000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 622) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000111111111110000000000000000111111111111100000000000000111111111111110000000000000111110000111111000000000000011110000000111000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111111000010000000000000000011111111111100000000000000000111111111110000000000000000001111111111000000000000000000111111110000000000000000000011111000000000000000000000001111000001110000000000000000111111111111100000000000000011111111111110000000000000000111111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 623) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000000111110000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000001111100000000000000000000001111100000000000000000000011111100000000000000000000001111100000000000000000000011111100000000000000000000011111100000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000000110000001111110000000000000011111111111111100000000000001111111111111100000000000000001111100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 624) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111111111000000000000001111111111111110000000000001111111111111111100000000001111110000011111110000000000111100000000111111000000000011100000000001111100000000001111000000000001100000000000111111111100000000000000000001111111111000000000000000000011111111110000000000000000001111111110000000000000000001111111000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000000011111111100000000000000000001111111110000000000000000000111111111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 625) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000011111100000000000000000000111111000000000000000000000111111000000000000000000000011111100000000000000000000011111100000000000000000000001111100000000000000000000000111100000000000000000000000011110000000110000000000000001111111111111110000000000000111111111111111000000000000001111111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 626) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111100000000000000000111111111110000000000000000011111111111000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000011111000000000000000000000001111111000000000000000000001111111100000000000000000001111111110000000000000000000111111110000000000000000000111110000000000000000000000011111000000000000000000000000111111100000000000000000000011111111000000000000000000000111111100000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 627) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000111110000000000000000000000111111000000000000000000000111111000000000000000000000111111000000000000000000000011111000000000000000000000011111100000000000000000000001111100000000000000000000001111100000000000000000000000111110000000000000000000000111110000000000000000000000111111000000000000000000000011111000000000000000000000001111000000000000000000000011111100000000000000000000011111110110000000000000000011111111111110000000000000000111111111111000000000000000011111111111100000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 628) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000111111111110000000000000000111111111111000000000000000111111100000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111111000000000000000000000001111111111000000000000000000011111111100000000000000000000111111110000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011111111100000000000000000001111111110000000000000000000011111111000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 629) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000111000000000000000001111111111110000000000000001111111111111000000000000001111111111111000000000000000111111100000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 630) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000111111111100000000000000000111111111110000000000000000011111111111000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111111100000000000000000000111111111000000000000000000011111111100000000000000000000111111000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011111111111000000000000000000111111111100000000000000000011111111111000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 631) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000111111110000000000000000000111111111100000000000000001111111111110000000000000000111111100100000000000000000111110000000000000000000000111110000000000000000000000011110000000000000000000000000111111111000000000000000000011111111100000000000000000000111111110000000000000000000011111111000000000000000000011111110000000000000000000001111100000000000000000000001111100000000000000000000000111111111111000000000000000011111111111100000000000000000111111111110000000000000000001111111111000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 632) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000001111100000000000000000000001111100000000000000000000000111111110000000000000000000111111111100000000000000000011111111110000000000000000001111111111000000000000000000011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 633) begin
            pixels = 784'b0000000000000000000000000000000000000000000100000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011111111100000000000000000011111111110000000000000000001111111111000000000000000000111111111000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 634) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000011111111110000000000000000111111111111100000000000000111111111111110000000000000011111111111110000000000000011111111111110000000000000001111100000000000000000000001111110000001000000000000000111111111111110000000000000011111111111111100000000000000111111111111110000000000000011111111111110000000000000000111111111111000000000000000001111111111100000000000000000111111111111100000000000000011111111111110000000000000001111111111111000000000000000011111111111100000000000000001111111111000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 635) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001110000000000000000000111111111110000000000000000011111011111000000000000000011110000001100000000000000001110000000000000000000000000110000000000000100000000000001100000000000000000000000000111000111000000000000000000011111111100000000000000000001111111110000000000000000011111100000000000000000000011111000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111111111111100000000000000000111111111111000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 636) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000011100000000000001110000000001110000000000001111111001111111000000000000011111111111111000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 637) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000111111000000000000000000001111111100000000000000000011110000110000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000100000000000000000011111111110000000000000000000111111111000000000000000000011111000000000000000000000011110000000000000000000000011110000000000000000000000011100000000000000000000000001111000000000000000000000000111111111100000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 638) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000100000000000000000011111111111110000000000000001111111111111000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 639) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000001111111111111100000000000011111111111111111000000000111110000000001111100000000011100000000000011100000000001110000000000000010000000000111000000000000000000000000011100000000000000000000000000111000111110000000000000000001111111111100000000000000000111111111110000000000000000011111111111000000000000000111111111110000000000000000111100000000000000000000000011110000000000000000000000001111111000000111100000000000011111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 640) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000001000000000000000111000000011110000000000000011111111111100000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 641) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000111000000000000000001111111111000000000000000001111111111000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 642) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000111111111000000000000000001111111111100000000000000011111000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000001111111111000000000000000000111111111000000000000000000111111111100000000000000000111110000000000000000000000111110000000000000000000000011100000000000000000000000001111111111100000000000000000111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 643) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111111110000000000000000001111111111100000000000000001111100111110000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000011000000000000000000000000001111111111100000000000000000111111111111000000000000001111111111111100000000000000111111111111100000000000000111110000000000000000000000111100000000000000000000000111100000000110000000000000001111111111111110000000000000111111111111111000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 644) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000001111111111111110000000000001111110000001111000000000001111100000000000000000000001111000000000000000000000000111000000000000000000000000011100000000100000000000000000111000011111000000000000000011111111111100000000000000000111111111100000000000000000011111100000000000000000000011111000000000000000000000111110000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000000111110000000000000000000000001111111111111111100000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 645) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111000000000000000000111111111100000000000000000111100001111000000000000000111100000001000000000000000111100000000000000000000000011100000000000000000000000001100000000000000000000000000111000000000000000000000000011110001110000000000000000000111111111100000000000000000001111111100000000000000000000011111100000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000011110000000010000000000000001111111111111100000000000000011111111111100000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 646) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000011111111000000000000000001111111111110000000000000001111110000111110000000000001111000000001111000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000001110000011110000000000000000111111111111000000000000000001111111111100000000000000000111111111100000000000000000011111000000000000000000000011110000000000000000000000001110011110000000000000000001111111111100000000000000000111111111100000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 647) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000011100100000000000000111111111111111000000000000111111111111111000000000000011111000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 648) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000010000000000000000111000000011100000000000000011111110111100000000000000001111111111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 649) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000111111110000000000000000001111111111100000000000000011111000001110000000000000011111000000011000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011110000000000000000000000001111110000000000000000000000011111111100000000000000000011111111110000000000000000111111000011000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000011110001111111111100000000001111111111111111110000000000011111111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 650) begin
            pixels = 784'b0000000000000000000000000000000000000000000111100000000000000000000000111110000000000000000000000011111000000000000000000000011111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000111110000000000000000000000011110000000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000110000000000000111000000000111000000000000111100000000011100000000000011110000011111110000000000001111111111111110000000000000011111111111110000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 651) begin
            pixels = 784'b0000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000010000000000000000111000111111111000000000000011111111111111000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 652) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000111111111100000000000000001111111111111000000000000001111000000111000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011110000000000000000000000011111111110000000000000000111111111110000000000000000111110000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000111111111100000000000000000000111111111000000000000000000000001111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 653) begin
            pixels = 784'b0000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011000000001110000000000000001100000001110000000000000001100000001100000000000000000110000001100000000000000000011111111100000000000000000001000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 654) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000001100000000000001110000000001110000000000001110000000001110000000000000110000000001110000000000000011111111111110000000000000001111111111110000000000000000000110111100000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 655) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111110000000000000000000011111111110000000000000000011110000111110000000000000011110000001111100000000000011110000000001110000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111100111100000000000000000001111111110000000000000000000111111111000000000000000000011111111100000000000000000011111000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111111111111111100000000000001111111111111110000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 656) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000111111111000000000000000000111111111110000000000000000111100000111100000000000000111100000011110000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001111011100000000000000000000011111111000000000000000000001111111110000000000000000000111111110000000000000000000111100110000000000000000000111100000000000000000000000111100000000000000000000000011111111000000000000000000000111111111110000000000000000000000011111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 657) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000010000000000000000011000000011000000000000000011000000011100000000000000001111000011000000000000000000011111111100000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 658) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000011111100000000000000000000111111111000000000000000000111100011100000000000000001111000001111000000000000000111000000111100000000000000111000000000111000000000000011000000000000000000000000001100000000000000000000000000111101111111000000000000000001111111111110000000000000000111111111110000000000000000011111000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000011100000000000000000000000001111110000011000000000000000011111111111110000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 659) begin
            pixels = 784'b0000000000000000000000000000000000000000000000100000000000000000000000000110000000000000000000000000111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000011000000000000001110000000111100000000000000111111100111000000000000000000111111111000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 660) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000011111111100000000000000001111111111110000000000000001111111110110000000000000000111110000000000000000000000111110000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100001111111000000000000001111111111111100000000000000011111111111111111110000000000111111111111111111000000000011111111111111111100000000011111111111111111000000000001111111111111110000000000000111110011111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 661) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000111100000000000000000000000011111000000000000000000000011111100000000000000000000001111100000000000000000000001111100000000000000000000000111100000000000000000000000111110000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000000111110001111101100000000000011111111111111111100000000000111111111111111110000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 662) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000111111111100000000000000011111111111100000000000000111111111100000000000000011111111100000000000000000011111100000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000001111111000000000000000000000111111111110000000000000000000111111111100000000000000000000111111110001111000000000001111111111111111100000000001111111111111111100000000001111111111111111100000000000111111111111100000000000000000111111111000000000000000000011111110000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 663) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000011111000000000000000000000111111000000000000000000000110111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001111100000000000000000000000111111111111110000000000000000111111111111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 664) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000001111111111111000000000000001111111111111000000000000001111100000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100011000000000000000000000111111100000000000000000000011111110000000000000000000001111000000011100000000000001111000011111110000000000001111000111111110000000000000111111111111100000000000000001111111111000000000000000000000111110000000000000000000000011110000000000000000000000001110000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 665) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000111111000000000000000000000011111100000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111110000000000000000000000001111111100000000000000000000000111111110000000000000000000000000111111000000000000000000000001111110000000000000000000000011111000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 666) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000011111111111000000000000001111111101111000000000000000111111000000000000000000000111110000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001111110001100000000000000000011111111110000000000000000000011111111000000000000000000011111110000000000000000000111111000000000000000000000011110001111111000000000000111111111111111100000000000011111111111111000000000000001111111111100000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 667) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000111111111111100000000000000011111111111110000000000000001100000000000000000000000000111100000000000000000000000001111000000000000000000000000011110000000000000000000000000011110000000000000000000000000111111100000000000000000000000111111000000000000000000000001111100000000000000000000000111110000000000000000000001111110000000000000000000011111100000111000000000000001111011111111110000000000001111111111111100000000000001111111111111000000000000000111111111100000000000000000001111111000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 668) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000011111111111100000000000000011111000000110000000000000011110000000010000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001111000000001000000000000000011111001111100000000000000000011111111110000000000000000000111111100011000000000000000111110011111110000000000000111111111111110000000000000011111111111000000000000000011111111110000000000000000000111111110000000000000000000001111100000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 669) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000111100000000000000000000011111110000000000000000000011111110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111110000000000000000000000111111111111110000000000000001111111111111110000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 670) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001111100000000000000000000011111100000000000000000000111111000000000000000000000011111000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001111111111000000000000000000011111111111111111000000000000000000111111111111000000000000000000011111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 671) begin
            pixels = 784'b0000000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000110011000000000000000111111111001100000000000000001111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 672) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000011111111111111000000000000111111110000011100000000000111110000000001100000000000111100000000001100000000000011100000000001000000000000001110000000000000000000000000011100000000000000000000000001111000000000000000000000000011110000000000000000000000000111111111000000000000000000000111111100001100000000000000011111000111110000000000000001110001111110000000000000001111111111100000000000000001111111111100000000000000000111111111100000000000000000000011110000000000000000000000001111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 673) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000001111111111000000000000000011111100001100000000000000001110000001100000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011000001111000000000000000000111111111100000000000000000001111100000000000000000000001111000000000000000000000001111000001111110000000000000111001111111110000000000000011111111111000000000000000001111111111000000000000000000000011110000000000000000000000011100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 674) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000001111111111000000000000000001111110111100000000000000011110000011100000000000000011100000011100000000000000001100000000000000000000000000111000000000000000000000000001110000000000000000000000000011110000000000000000000000000111111110000000000000000000000111111000000000000000000000111100000000000000000000000111000000111100000000000001111111111111110000000000001111111111111000000000000000111111111110000000000000000000000111100000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 675) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000001111100000000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111111111101000000000000000011111111111111111100000000000111111111111111111000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 676) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111100000000000000000000011111110000000000000000000011111100000000000000000000011111100000000000000000000011111000000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001111000000000000000000000000111110000000000000000000000001111111111111000000000000000011111111111111110000000000000000111111111111100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 677) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111000000000000000001111110111000000000000000011111000000000000000000000011110000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001110000000000000000000000000111101000000000000000000000000111111111100000000000000000000001111100000000000000000000001111000000000000000000000001111101111100000000000000001111111111110000000000000001111111111110000000000000000111111111100000000000000000000011111100000000000000000000001110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 678) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000011110000000000000000000000000111000000000000000000000000011100000000000000000000000111110000000000000000000000011110000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111111110000000000000000000001111111111110000000000000000000111111111100000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 679) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000011111111100000000000000001111111111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000011111100000000000000000000001111000000000000000000000011111000000000000000000000001111000000000000000000000000111000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001111111100000000000000000000011111111110000000000000000000001111111111100000000000000000001111111111000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 680) begin
            pixels = 784'b0000000000000000000000000000000000000000000011110000000000000000000000011110000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000011111100000000000000000000000111111111111111110000000000000111111111111111000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 681) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000011111111111110000000000000011111000000011100000000000011100000000000111000000000011100000000000011100000000001110000000000000110000000000111000000000000000000000000001110000000000000000000000000011000000000000000000000000000110000000000000000000000000001111111100000000000000000000111111100000000000000000000001111000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111111111100000000000000000001111111110000000000000000000011111111000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 682) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000111111111111000000000000001111110000111111000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011111111111111000000000000000111111111111100000000000000000000111111000000000000000000000011110000000000000000000000111110000010000000000000000111111111111111100000000000011111111111111110000000000000100000111111100000000000000000011111110000000000000000000011111000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 683) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000111111110000000000000000000111111111100000000000000000011110001110000000000000000011110000110000000000000000011110000010000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011110000000000000000000000001111100011100000000000000000011111111110000000000000000001111111111000000000000000000111111111100000000000000000011111100000000000000000000011110000000000000000000000001110000000000000000000000000111111111111100000000000000011111111111110000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 684) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000001100000000000000011100000001110000000000000011100000001110000000000000011110000001111000000000000001111011111111100000000000001111111111111100000000000000011111111111100000000000000001111000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 685) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000011111111100000000000000000111111111111000000000000000111111111111100000000000000011111000001110000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000001111000000000000000000000000111110000000000000000000000011111111000000000000000000000111111111111000000000000000001111111111100000000000000000001111111100000000000000000000111111000000000000000000000111111111111000000000000000011111111111100000000000000001111111111110000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 686) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000111000000000001111000000000111110000000000111100000000111110000000000111100000001111110000000000011100000111111110000000000001111111111111110000000000000111111111111110000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 687) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111110000000000000001111111111111100000000000000111110000001111000000000000111100000000011100000000000111000000000000110000000000111100000000000011000000000011110000000000000000000000001111000000000000000000000000011100000000000000000000000001111100000111100000000000000011111111111111000000000000000111111111111100000000000000011111111111100000000000000001111111100000000000000000001111100000000000000000000000111111110000000000000000000011111111000000000000000000001111111100000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 688) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111111111111100000000000000011111111111110000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 689) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001111111111111100000000000001111110000111110000000000001111000000000011000000000001110000000000011100000000000111000000000001100000000000111000000000000000000000000001110000000000000000000000000111000000000000000000000000001110000000000000000000000000111111111100000000000000000001111111111000000000000000000011111111000000000000000000011111000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000011111111110000000000000000001111111111000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 690) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000010000000000000001111100000111000000000000000111110000111100000000000000111111111111100000000000000011111111111100000000000000001111111111110000000000000000111111111110000000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 691) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000001111111000000000000000000001111111110000000000000000001110000011000000000000000001110000001100000000000000000110000000100000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011100000111110000000000000001111111111111000000000000000011111111111000000000000000001111111100000000000000000000111110000000000000000000000111100000000000000000000000011100000000000000000000000011000000111100000000000000001110111111110000000000000000111111111100000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 692) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000011111000000000000000000000011111100000000000000000000011111100000000000000000000011011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000011000000000000001111000000011100000000000001111100000111110000000000000111000000111111000000000000011000000011111000000000000011100011111110000000000000011111111111110000000000000001111111111110000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 693) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000001111110000000000000000000001100110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000001000000000000001100000000001110000000000001110000000001110000000000000110000000001110000000000000110000011111111000000000000111011111111111100000000000111111111111111100000000000011111111110101100000000000011110000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 694) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000011111111000000000000000000011111001100000000000000000111100000110000000000000000111100000111000000000000000011100000011000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000001111000000000000000001111111111100000000000000000111111111100000000000000000001111111000000000000000000000111100000000000000000000000011100000000000000000000000011100000001000000000000000001110000001110000000000000000111000111111000000000000000011111111111000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 695) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000001111111111110000000000000001111100000011100000000000001110000000000011000000000001110000000000000110000000001110000000000000001000000001110000000000000001100000000110000000000000000110000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000001110000000000000000000000000111111111111100000000000000001111111111100000000000000000001111111000000000000000000000111000000000000000000000000011101111000000000000000000001111111110000000000000000000011111111000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 696) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000111100000000000000000000000111110000000000000000000000110110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000010000000000000001100000000011000000000000001110001011111100000000000000111111111111110000000000000011111111111110000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 697) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001000000000000100000000000000100000111111111000000000000011111111111111100000000000001111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 698) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000011111100000000000000000000001111110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000001110000000000000111000000000111000000000000111000000000111100000000000011000000100111100000000000011111111111111100000000000011111111111111110000000000000111100000111110000000000000000000000000111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 699) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000001111100000000000000000000000111110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000001110000000000001110000000001110000000000000111000000011111000000000000111000001111111000000000000011111111111111000000000000001111111111111000000000000000111111110010000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 700) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000001111111111111000000000000001111111111111111000000000001111100000000111100000000000111000000000000111000000000111000000000000011000000000011100000000000000100000000001110000000000000000000000000111100000000000000000000000001111000000000000000000000000011111100000000000000000000000111111111110000000000000000001111111111000000000000000000111111111100000000000000000111110000000000000000000000111100000000000000000000000011100000011100000000000000001111111111111000000000000000111111111111100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 701) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000001111111111000000000000000001111110011110000000000000000111000000011000000000000000111000000001100000000000000011100000001110000000000000011100000000110000000000000001110000000000000000000000000110000000000000000000000000011100000111000000000000000001111111111100000000000000000011111111110000000000000000001111111110000000000000000000111111000000000000000000000011100000000000000000000000001110000000000000000000000001100000011100000000000000000111111111110000000000000000011111111111000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 702) begin
            pixels = 784'b0000000000000100000000000000000000000001111000000000000000000000001111100000000000000000000000111110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000110000000000011100000000000111000000000011100000000000011000000000011100000000000011100000000001110000011111111110000000001111111111111111110000000000111111111111111111000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 703) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000011111111100000000000000000011111001111000000000000000001110000001100000000000000000110000000110000000000000000011000000001000000000000000011100000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000011100000000000000000000000001111111000000000000000000000001111111111000000000000000000011111111100000000000000000001111110000000000000000000001111000000000000000000000001111000001110000000000000000111101111111100000000000000001111111111100000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 704) begin
            pixels = 784'b0000000000000000000000000000000000000000111100000000000000000000000111110000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000011000000000000111111111111111110000000000011111111111111111000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 705) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000001111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000011000000000000011110000000011110000000000001110000000011110000000000001110000000001111000000000000110000000001111000000000000111000000001111100000000000111100001111111100000000000011111111111111100000000000011111111111111110000000000000111000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 706) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111110000000000000000111110000011000000000000000111100000000110000000000000011100000000010000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000001111111000000000000000000000011111111000000000000000000011111111100000000000000000011110000000000000000000000011100000000000000000000000011100000100000000000000000001110001111000000000000000000011111111100000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 707) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000011111111111100000000000000011111100011111000000000000011110000000011100000000000011110000000000111000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000111100000000000000011111111111110000000000000000111111111110000000000000000001111111110000000000000000000111111000000000000000000000111000000111000000000000000111000000011100000000000000011100000111110000000000000001101111111110000000000000000111111111000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 708) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000111111111110000000000000000111100000111110000000000001110000000000011110000000001110000000000000001100000000110000000000000000000000000011100000000000000000000000000111100000000000000000000000001111111111000000000000000000001111111100000000000000000000111100000000000000000000000011100000010000000000000000011111111111100000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 709) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000111111110000000000000000001111001111100000000000000000111000001110000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011110000000000000000000000000111100000000000000000000000000111110000000000000000000000011111000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000011000000000000000001110000011100000000000000000011111111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 710) begin
            pixels = 784'b0000000000000000000000000000000000000000111000000000000000000000000111110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000110000000000111111111111111111000000000000111111111111111100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 711) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111111100000000000000000011111111110000000000000000011110000111000000000000000001110000011100000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011110000000000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000001110000000000000000001111111111000000000000000000111111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 712) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001111110000000000000000000000111111000000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000001111000000000000000000000001111100000000000000000000000111111111100000000000000000011111111111111000000000000001111111111111110000000000000011111111111111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 713) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111100000000000000001111111111110000000000000001111000001110000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000001110111100000000000000000000111111111000000000000000000001111111100000000000000000001111111100000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000001110000110000000000000000000111111111000000000000000000001111111100000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 714) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000111110000000000000000000000011111100000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000001111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000001111100000000000000000000000111110000000000000000000000111111000000011000000000000011111111111111110000000000001111111111111111000000000000111111111111111000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 715) begin
            pixels = 784'b0000000000000000000000000000000000000000111000000000000000000000000111110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111110000000000000000000000111111100000000000000000000111111111111111100000000000011111111111111111100000000000111111111111111110000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 716) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000011111111100000000000000000011111111111000000000000000001111000111110000000000000001111000001111100000000000000111100000011100000000000000011110000000000000000000000000111000000000000000000000000011110000000000000000000000000111111100000000000000000000011111111000000000000000000001111111000000000000000000000111111100000000000000000000011100000000000000000000000011100000000000000000000000000110000000000000000000000000011100000000000000000000000000111111111110000000000000000011111111110000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 717) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000011111110000000000000000000011111111100000000000000000011111111111000000000000000001111101111100000000000000000111100011110000000000000000011100000111000000000000000001110000000000000000000000000111100000000000000000000000011111111100000000000000000001111111110000000000000000000011111111000000000000000000000111111000000000000000000000011110000000000000000000000001111000000000000000000000000111100001100000000000000000011111111111000000000000000001111111111100000000000000000011111111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 718) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001111111100000000000000000001111111111000000000000000000111111111110000000000000000011100111111100000000000000001110000111111000000000000000111000000111000000000000000111100000001000000000000000001110000000000000000000000000111101100000000000000000000011111111000000000000000000000111111100000000000000000000011111100000000000000000000001111100000000000000000000001111000000000000000000000000111100000000000000000000000011110001110000000000000000001111111111100000000000000000011111111110000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 719) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111100000000000000000000111111111000000000000000000111111111110000000000000000011110001100000000000000000011111000000000000000000000001111000000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000001111111000000000000000000000011111100000000000000000000011111110000000000000000000011111111000000000000000000000111110000000000000000000000011110000000000000000000000001111001110000000000000000000111111111100000000000000000001111111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 720) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000001111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000001111100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000011111000000000000000000000011111111111100000000000000001111111111111000000000000000011111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 721) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111100000000000000000111111111111000000000000000111100001111110000000000000111100000011111000000000000011110000001111100000000000011111000000111110000000000001111000000011110000000000000111110000000000000000000000011111000000000000000000000000111110000000000000000000000011111100000000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000000000000001111111110000000000000000000111111111000000000000000000011111110000000000000000000001111100000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 722) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011111000000000000000000000011111100000000000000000000001111110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000000111100000000000000000000000011110000000000000000000000001111111111000000000000000000111111111110000000000000000011111111111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 723) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011111111111111110000000000000111111111111110000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 724) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111111100000000000000001111111111111000000000000000111110011111100000000000000111110000111110000000000000011110000001110000000000000011111000000000000000000000001111100000000000000000000000111110011000000000000000000001111111111000000000000000000111111111000000000000000000001111111100000000000000000000111111000000000000000000000011111000000000000000000000001111100000000000000000000000111110000001000000000000000011111000001111000000000000001111111111111100000000000000111111111111100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 725) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000000111100000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000001111100000000000000000000000111110000000000000000000000111111000000000000000000000011111000001100000000000000001111110011111100000000000000111111111111110000000000000011111111111110000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 726) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111110000000000000000000000001111100000000000000000000000111111111100000000000000000000111111111000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 727) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111110000000000000000000111111111100000000000000000011100001110000000000000000011000000011100000000000000001100000000110000000000000000110000000011000000000000000011000000000000000000000000001110000000000000000000000000011100000000000000000000000001111000000000000000000000000111110000000000000000000000111111000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000001100000000000000000000000000111111110000000000000000000001111111000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 728) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000111110000000000000000000000011110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000001111111100000000000000000000111111111110000000000000000011111111111000000000000000000111111111100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 729) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000001111111111111110000000000001111111111111111100000000000111000000000011110000000000011100000000000110000000000011110000000000000000000000001110000000000000000000000000011100000000000000000000000000111000000000000000000000000011111000000000000000000000000111110000111000000000000000000011111111110000000000000000001111111110000000000000000011111100000000000000000000011111000000000000000000000001111000000000000000000000000011110000000110000000000000001111111111111000000000000000011111111111000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 730) begin
            pixels = 784'b0000000000000000000000000000000000000011110000000000000000000000001111000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000001100000000000001100000000000110000000000000111001110001111000000000000111111111111111100000000000011111111111111100000000000000110000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 731) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000011111100000011110000000000011111000000000011000000000001110000000000000110000000000111000000000000001000000000011100000000000000100000000001110000000000000010000000000111000000000000000000000000011110000000000000000000000000111100000000000000000000000001111100000000000000000000000001111111111000000000000000000111111111100000000000000000111111110000000000000000001111100000000000000000000000111000001111000000000000000111111111111111100000000000011111111111111111000000000000111100000000111100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 732) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011111111111000000000000000001111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 733) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000011111100000111000000000000001110000000000110000000000001100000000000011100000000001110000000000000111000000000110000000000000001100000000011000000000000000110000000001100000000000000000000000000110000000000000000000000000001100000000000000000000000000111000000000000000000000000001110000111110000000000000000011111111110000000000000000000111111100000000000000000001111110000000000110000000001111000000000001111000000000111000000000001111000000000001110000000111111000000000000111111111111100000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 734) begin
            pixels = 784'b0000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000001100000000011000000000000001110000000001110000000000001111000000000111111111111111111000000000010111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 735) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111111100000000000000000011110000111000000000000000011100000000110000000000000001100000000001100000000000000111000000000110000000000000011100000000011000000000000000110000000011100000000000000011100000000000000000000000000111000000000000000000000000011110000000000000000000000000011111110000000000000000000001111111000000000000000000001111100000000000000000000011111000000000000000000000001110000000000000000000000000111000000000000000000000000011100000111000000000000000001111111111000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 736) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000001100000000000000000110000011111000000000000000111111111111000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 737) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000011111111100000000000000000011100000111000000000000000011100000000110000000000000001110000000011000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011100111000000000000000000000111000000000000000000000000011111111100000000000000000001111111100000000000000000001111000000000000000000000001110000000000000000000000000110000000000000000000000000111000000011100000000000000011000000011110000000000000000110000011110000000000000000011111111110000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 738) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111110000000000000000011110000011100000000000000001100000000110000000000000000110000000001000000000000000011000000000100000000000000001100000000110000000000000000110000000000000000000000000011100000000000000000000000001111111111110000000000000000111111111111000000000000000000111111110000000000000000000111110000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000011000000111000000000000000001110001111100000000000000000011111111000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 739) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111110000000000000000111110000111110000000000000111000000000011100000000000011000000000000111000000000001100000000000001100000000000110000000000000110000000000011000000000011110000000000001100000000000000000000000000011000000000000000000000000000110011111100000000000000000001111111111000000000000000000111111110000000000000000001111110000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011100000001110000000000000000111111111111000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 740) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000001110000000000000000000000000111000000000000000000000000011111111100000000000000000000111111111100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 741) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000011111111100000000000000000011100001111000000000000000011100000001100000000000000001100000000010000000000000000110000000011000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000011000000000000000000000000001111111110000000000000000000111111111100000000000000000111111111100000000000000000011000000000000000000000000001100000001100000000000000000110000111110000000000000000011111111110000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 742) begin
            pixels = 784'b0000000000000000000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000000111000000000000000000000000011100000000001100000000000000110000001111110000000000000011111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 743) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000011100000000000001100000000011110000000000001110000000111100000000000000111000000111100000000000000011100001111000000000000000000111111110000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 744) begin
            pixels = 784'b0000000000000000000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000111000000000000001110000001111100000000000000011000011111110000000000000001111111011100000000000000000001110001100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 745) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000011111111111100000000000000011110000000111000000000000011100000000011100000000000001100000000001110000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001110000000000000000000000000011000000000000000000000000001110000000000000000000000000011100000110000000000000000000011111111100000000000000000011111100000000000000000000011110000000000000000000000001100000000110000000000000000110000000011000000000000000011100001111000000000000000000111111111000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 746) begin
            pixels = 784'b0000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000110000000000000110000000011111000000000000001100000111110000000000000000111111111110000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 747) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000001000000000000011100000000111100000000000001100000000111110000000000001110000001111100000000000000111111111111000000000000000011111111100000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 748) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000001000000000000110000000000001110000000000111000011111111110000000000011111111111111100000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 749) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000011100000000000011100000000011110000000000001110000000011110000000000000110000001111110000000000000011000111111110000000000000001111111100000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 750) begin
            pixels = 784'b0000000000000000000000000000000000000000000100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000001100000000000000110000000011110000000000000011000000111110000000000000001111111111110000000000000000001111000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 751) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000011111111111000000000000000111110000000110000000000000111100000000001100000000000011100000000000010000000000001100000000000001000000000000110000000000000100000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000001100000000000000000000000000011001111110000000000000000000111111111000000000000000000001110010000000000000000000001110000000000000000000000000110000000001100000000000000011000000001100000000000000001110000111100000000000000000011111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 752) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111111000000000000000111100000111110000000000000111000000000111000000000000011000000000000000000000000011100000000000000000000000000110000000000000000000000000111000000000000000000000000001100000000000000000000000000111000000000000000000000000001110011111000000000000000000011111111100000000000000000001111111000000000000000000000111000000000000000000000000111000000000000000000000000011100000000110000000000000001100000111111000000000000000111111111111000000000000000001111111100000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 753) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000111111100000000000000000000111111111100000000000000000111111111110000000000000000111100000111000000000000000011100000011100000000000000001110000001100000000000000000110000000000000000000000000011100000000000000000000000001111001110000000000000000000111111111000000000000000000001111111100000000000000000000011111110000000000000000000001111100000000000000000000000111000000000000000000000000011000000000000000000000000001111111100000000000000000000111111110000000000000000000011111111000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 754) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000010000000000000000111000000111100000000000000011100001111110000000000000001110111111110000000000000001111111111110000000000000000111111111110000000000000000001110000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 755) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000001111111110000000000000000001111111111110000000000000000111111111111100000000000000011100001111110000000000000001110000000111000000000000000111000000001000000000000000011111000000000000000000000000111111110000000000000000000011111111000000000000000000001111111100000000000000000001111111100000000000000000001111100000000000000000000001111100000000000000000000000111000000000000000000000000011100001100000000000000000001111111110000000000000000000111111111000000000000000000001111111000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 756) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000110000000000000000011111111111100000000000000001111111111110000000000000000011111111110000000000000000000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 757) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111000000000000000001111111111100000000000000001111111111110000000000000000111100000011000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011111110000000000000000000001111111100000000000000000000011111110000000000000000000000111110000000000000000000000111110000000000000000000000011100000010000000000000000001110000111100000000000000000111111111110000000000000000011111111110000000000000000000111111110000000000000000000011111110000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 758) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000111110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000001100000000000000111000000011110000000000000111100000011111000000000000011100001111111000000000000001111111111111000000000000001111111111110000000000000000111111110010000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 759) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000011111111000000000000000000111111111110000000000000000011110000110000000000000000011100000011000000000000000011100000001000000000000000001110000000000000000000000001111000000000000000000000000011110000110000000000000000001111111111000000000000000000011111111100000000000000000000011111100000000000000000000011111000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000000111000001110000000000000000011111111111000000000000000000111111111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 760) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111100000000000000000111111111111000000000000001111100000111100000000000001111000000001100000000000000111000000001110000000000000111100000000110000000000000011110000000000000000000000001111000000000000000000000000011111000000000000000000000000111111110000000000000000000001111110000000000000000000000011111000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011110000000000000000000000001111111110000000000000000000011111111000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 761) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000111111111100000000000000001111111111110000000000000001111110000111000000000000000111100000011100000000000000111100000001100000000000000011110000000000000000000000000111100000000000000000000000011111111110000000000000000000111111111000000000000000000000111111000000000000000000000011111000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011111011110000000000000000000111111111000000000000000000001111111000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 762) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000001111111100000000000000000001111111111000000000000000001111111111100000000000000000111000011100000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011111000111100000000000000000111111111100000000000000000001111111100000000000000000000001111100000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001111000000000000000000000000011111111000000000000000000001111111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 763) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111111000000000000000111111111111100000000000000011111110111110000000000000011110000000110000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000001111011111000000000000000000111111111110000000000000000011111111100000000000000000000111111110000000000000000000011111000000000000000000000011100000000000000000000000011110000000000000000000000000111000000000000000000000000011111111111000000000000000001111111111000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 764) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001110000000001100000000000001111000001111110000000000000111111111111111000000000000111111111111110000000000000011111111111110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 765) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000111000000000000000110000000011100000000000000011000111111100000000000000011111111111100000000000000001111111110000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 766) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000011100000000000001110000000111110000000000000110000111111110000000000000111001111111110000000000000011111111111000000000000000001111100000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 767) begin
            pixels = 784'b0000000000000000000000000000000000000000111100000000000000000000000111110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011111111111111110000000000001111111111111111000000000000011111111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 768) begin
            pixels = 784'b0000000000000000000000000000000000000000000111100000000000000000000000111110000000000000000000000111110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100001100000000000000000011110001110000000000000000011111111111100000000000000001111111111110000000000000000111111111110000000000000000011111111110000000000000000000111110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 769) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000111100000000000000000000001111110000000000000000000000111111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000001110000000000000001110000111111000000000000000111001111111100000000000000011111111111100000000000000001111111111000000000000000000111111110000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 770) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000111000000000000001111000001111100000000000000111001111111100000000000000011111111111100000000000000001111111111000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 771) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000001111111111000000000000000001111111111100000000000000011111111111110000000000000001111100000011000000000000001111100000001000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111110000000000000000000000011111100000000000000000000001111110000000000000000000000111111000000000000000000000111110000000000000000000000011110000000000000000000000001110000000000000000000000000111100010000000000000000000011111111100000000000000000000111111100000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 772) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000111111111110000000000000000011111111111100000000000000011111000001111000000000000011100000000001100000000000001110000000000100000000000000110000000000000000000000000011000000000000000000000000001110000110000000000000000000011111111100000000000000000001111111100000000000000000000011111110000000000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000001110000000000000000000000000111111111000000000000000000001111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 773) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000111110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000001100000000000000111000000011111000000000000011100001111111000000000000001111111111111000000000000000111111111111000000000000000011111011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 774) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111111000000000000000011111111111000000000000000001111111000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011110011110000000000000000000111111111000000000000000000011111111000000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000000111000001100000000000000000011111111111100000000000000001111111111100000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 775) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111100000000000000000111111111111000000000000000011111101111100000000000000011110000000100000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000011111110000000000000000000000111111100000000000000000000001111110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000001100000000000000001111111111111000000000000000011111111111100000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 776) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000001111111110000000000000000001111111111100000000000000001111111111110000000000000001111100000011000000000000001111100000001100000000000000111100000000100000000000000011100000000000000000000000001110000000000000000000000000111111110000000000000000000001111111100000000000000000000111111110000000000000000000011111110000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000001111110000000000000000000000111111000000000000000000000011111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 777) begin
            pixels = 784'b0000000000000000000000000000000000000000111100000000000000000000000111110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000011110000000000000001111111111111111000000000000111111111111111100000000000011111111111111110000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 778) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001111100000001000000000000000111111111111110000000000000001111111111111000000000000000011111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 779) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000001111111111111000000000000001111111111111100000000000001111100000000100000000000000111000000000000000000000000111100000000000000000000000001110000000000000000000000000111100000000000000000000000001111000000000000000000000000011110000000000000000000000000111111100000000000000000000011111110000000000000000000011111110000000000000000000011111000000000000000000000111110000000000000000000000011110000000000000000000000001110000011100000000000000000111111111110000000000000000011111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 780) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000011000000000000000011100111111100000000000000001111111111000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 781) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111110000000000000001111110011111100000000000001111000000001110000000000000111000000000011000000000000011000000000000000000000000001110000000000000000000000000111000000000000000000000000011110000000000000000000000000111100011000000000000000000001111111100000000000000000000001111100000000000000000000011111000000000000000000000011111000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011111000000000000000000000000111111110000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 782) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011111100000000000000000000000111111111110000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 783) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000001111111111111000000000000011111111111111100000000000011111100000000000000000000001111000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000001111000000000000000000000000111110000000000000000000000001111111111111000000000000000001111111111100000000000000000000111111110000000000000000000111111000000000000000000001111100000000000000000000001111100000000000000000000000111100000000000000000000000011111111111000000000000000000111111111110000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 784) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000110000000000000000011111111111000000000000000001111111111000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 785) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000100000000000000111000000001110000000000000111000000001111000000000000011100000011111100000000000011100000111111000000000000001110011111111000000000000000111111111000000000000000000011111110000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 786) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111100000000110000000000000011100000001111000000000000001110000001111000000000000000111000011111000000000000000011111111111000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 787) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111110000000000000000111111011111100000000000000011100000111110000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001110000000000000000000000000011110010000000000000000000000111111100000000000000000000011111100000000000000000000011111000000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001111000000011000000000000000011111111111100000000000000000111111111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 788) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111111110000000000000001111111111111100000000000001111100000001111000000000000111000000000011000000000000111100000000000000000000000001110000000000000000000000000111000000000000000000000000011110000000000000000000000001111000000000000000000000000011111001100000000000000000000111111111000000000000000000001111111000000000000000000001111100000000000000000000011111000000000000000000000011110000000000000000000000011110000011110000000000000001111111111111000000000000000011111111110000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 789) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000011111111111111000000000000011111111111111110000000000011110000000001110000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011100000000000000000000000001111000000000000000000000000011110101100000000000000000000111111110000000000000000000111111111000000000000000000111110000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111111101000000000000000000000111111111100000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 790) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000011111111111110000000000000001111111111111100000000000001111000000111110000000000000111000000001110000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000001110000000000000000000000000011100000000000000000000000001111111110000000000000000000011111111100000000000000000001111111110000000000000000011111110000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000000011111111111100000000000000001111111111110000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 791) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001111111111110000000000000001111110001111100000000000001111000000111110000000000000111000000000110000000000000011000000000000000000000000001110000000000000000000000000111000000000000000000000000001110000000000000000000000000111100000000000000000000000001111111100000000000000000000011111110000000000000000000001111111000000000000000000011111000000000000000000000011111000000000000000000000001110000000000000000000000000111000000000000000000000000011111111100000000000000000000111111110000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 792) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000011111111100000000000000000111111111110000000000000001111100000111000000000000000111000000111100000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001110000000000000000000000000011111111100000000000000000000111111100000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000000111111111000000000000000000011111111000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 793) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111111111000000000000001111111001111110000000000001111000000001111100000000001111000000011111110000000000111000000000111110000000000001110000000000000000000000000111000000000000000000000000011111000000000000000000000000111100001100000000000000000001111111111000000000000000000011111111100000000000000000001111111000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000001111000000000000000000000000111111110000000000000000000001111111000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 794) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000001110000000000001110000000011111000000000000111100001111111000000000000011111111111111000000000000000011111110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 795) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000111111000000000000111111111111111100000000000011111111111110000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 796) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000111111111110000000000000000111110011111100000000000000011100000001110000000000000011100000000111000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001110000000000000000000000000111100011000000000000000000001111111110000000000000000000011111110000000000000000000001111100000000000000000000001111000000000000000000000001111000000000000000000000001110000000000000000000000001111000000000000000000000000011111100000000000000000000001111111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 797) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001111111111111100000000000001111111111111111000000000001111100000000111110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 798) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000111100000000000000000000000011111111111000000000000000000111111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 799) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111111111111100000000000000001111111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 800) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111111000000000000000011111111111110000000000000001111000000111100000000000001111000000001100000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000001111000000000000000000000000011111111100000000000000000000111111110000000000000000000001111110000000000000000000001111100000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011111111110000000000000000000111111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 801) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000001110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000001110000000000011100000000001111000000000001110000000011111000000000001111000000111111000000000000111000001111111000000000000011111111111111000000000000000111111111111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 802) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000001111111111100000000000000001111111111111000000000000001111000000001110000000000000111000000000011000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111000001000000000000000000011111111110000000000000000000111111111000000000000000000011111100000000000000000000011111000000000000000000000011110000000000000000000000001111000000000000000000000000011111000000000000000000000000111111000000000000000000000000111110000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 803) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111111110000000000000000000011111111111100000000000000000111111111110000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 804) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000001111111100000000000000000111111111110000000000000000111110000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001110000011110000000000000000111111111110000000000000000001111111100000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000001110000000100000000000000000111000001110000000000000000011111111111000000000000000001111111111000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 805) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000010000000000000000111000000011100000000000000011000000011100000000000000011111111001110000000000000011111111111110000000000000001111000111110000000000000000100000001110000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 806) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000001111111110000000000000000011111100111000000000000000011110000000100000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000011000000000000000000011110111110000000000000000000111111110000000000000000000011111110000000000000000000000111000000000000000000000000111000000000000000000000000011000000110000000000000000011100011111000000000000000001110111111100000000000000000011111111110000000000000000000111111000000000000000000000011100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 807) begin
            pixels = 784'b0000000000000000000000000000000000000000000000010000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011111000000000000000000000011111000000001100000000000011111000000001110000000000011111000000001111000000000001111000000001111100000000001111111111011111000000000000111111111111111100000000000011111111111111110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 808) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000111100000000000000000000000011110000000111100000000000011110000000011100000000000011110000000111100000000000011110000000111100000000000011111111000111110000000000011111111111111100000000000000111111111111110000000000000000000000111100000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 809) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000111111111000000000000000000111100001110000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000001100001100000000000000000000111111110000000000000000000001111110000000000000000000000111100000000000000000000000011000000000000000000000000011100000000000000000000000011100000010000000000000000000110001111000000000000000000011111111100000000000000000000111111000000000000000000000111110000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 810) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000011111111111000000000000000111111111111111000000000000111100000000011100000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001110000001100000000000000000111111001110000000000000000001111111110000000000000000000011111100000000000000000000001111000000000000000000000001111000000000000000000000000111000111100000000000000000111111111110000000000000000011111111110000000000000000001111111000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 811) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000111111110000000000000000001111000000000000000000000000110000000000000000000000000011000000000000000000000000001000000000000000000000000001110000000000000000000000000111000000000000000000000000001100001100000000000000000000111111110000000000000000000011111110000000000000000000001111000000000000000000000001111100000000000000000000000111000010000000000000000000011100011100000000000000000001111111110000000000000000000011111100000000000000000000001111000000000000000000000011111000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 812) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000011100000000000000001111000001110000000000000001111111101110000000000000000111111111110000000000000000000000001110000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 813) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000111111111111000000000000011111111000111000000000000011111000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000010000000000000000001110000111100000000000000000111111111110000000000000000001111111100000000000000000000011111000000000000000000000001111000000000000000000000011110000000000000000000000011110000000000000000000000001110010111000000000000000000111000111100000000000000000011110111110000000000000000000111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 814) begin
            pixels = 784'b0000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000001000000000000000111100000011110000000000000111100000001111000000000000111110000001111000000000000111111110001111000000000000111111111111111000000000000001100000111110000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 815) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000011111111111110000000000000111111100000111000000000000111110000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000001000000000000000001111010011110000000000000000011111111110000000000000000001111111000000000000000000011111110000000000000000000111111100000000000000000000011110000000000000000000000011110000000000000000000000001110000000011100000000000000111111111111111000000000000001111111111111000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 816) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000001111111111111100000000000011111000000001110000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000011100000011000000000000000001111111111100000000000000000011111111100000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100001001100000000000000001111110111110000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 817) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000111100000000001000000000000011100000000001110000000000011100000000001111000000000011110000000001111000000000011111111110001111000000000011111111111111111000000000001100000001111111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 818) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000011111111111100000000000000111110000001111000000000000111000000000001100000000000111000000000001110000000000011000000000000110000000000011100000000000000000000000001110000000000000000000000000011000000100000000000000000001111111110000000000000000001111111110000000000000000001111100000000000000000000000111000000001100000000000000011000000111110000000000000011111111111110000000000000000111111111000000000000000000001111110000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 819) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111111111000000000000001100000000011110000000000001100000000000011000000000001110000000000000000000000000110000000000000000000000000011000001110000000000000000001100111111000000000000000000111111110000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000011100000011000000000000000001110000111110000000000000000011111111110000000000000000000001111000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 820) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000001000000011100000000000000000110000001100000000000000000011000001110000000000000000001100001110000000000000000000100001110000000000000000000010001110000000000000000000000001110000000000000000000000001110000000011100000000000000111000000011100000000000000111000000001110000000000000111100000001100000000000000011111111001110000000000000001111111111111000000000000000000000011111000000000000000000000000111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 821) begin
            pixels = 784'b0000000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011100000000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000110000000000001111000000000111000000000001111111111100111000000000000111111111111111100000000000000000000001111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 822) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000111111111111100000000000000111111100000000000000000000111110000000000000000000000011110000000000000000000000001111100000000000000000000000011111111100000000000000000000111111110000000000000000000001111111000000000000000000000011110000000000000000000000111110000000000000000000001111100000000000000000000001111100000000000000000000001111100000011110000000000001111000001111111000000000001111001111111111100000000001111111111111111000000000000111111111110000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 823) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000111100000000000000000000000011100111000000000000000000011111111100000000000011111111111111100000000001111111111111111100000000000111111111110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100111110000000000000000001111111111100000000000000000111111111110000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 824) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000111111111111111000000000000111110000000001000000000000111100000000000000000000000011100000000000000000000000001111000000000000000000000000011111111110000000000000000000011111111000000000000000000000011111100000000000000000000011111000000000000000000000111110000000000000000000001111100000000000000000000001111000000000000000000000001111000001111000000000000001111111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 825) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000001110000000000000000000000000111000000000000000000000000011101110000000000000000111111111111000000000011111111111111111000000000111111111011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011111111111000000000000000001111111111100000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 826) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000001110000000000000000000000001110000000000000000000000000011100100000000000000000000011100111000000000000000001111111111000000000011111111111111111100000000011111111111111110000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001110000000000000000000000001111000111111100000000000000111111111111110000000000000011111111111100000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 827) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000111111111111110000000000001111111110000010000000000011111100000000000000000000001110000000000000000000000000111000000000111000000000000001111111111111100000000000000111111111111110000000000000000000001111100000000000000000000001111000000000000000000000001111000000000000000000000011110000000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000111100000111100000000000000111111111111110000000000000011111111111110000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 828) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000110000000000000000000111011111100000000000000000111111111100000000000000011111111111000000000000001111111111000000000000000001111111100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000111100000000000000011101111111110000000000000001111111111100000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 829) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000001111111100000000000000000111111111000000000000000001111111000000000000000000001111100000000000000000000000111000000000000000000000000011000000000000000000000000001110000000000000000000000000111111110000000000000000000001111111000000000000000000000001111100000000000000000000011111000000000000000000000111110000000000000000000000111110000000000000000000001111100000000000000000000001111000000000000000000000001111000011110000000000000000111111111111000000000000000011111111111000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 830) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000100000000000000000001110111111000000000000000011111111111000000000000001111111111100000000000000011111111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011000001011000000000000000011111111111100000000000000001111111110000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 831) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110001100000000000000000000111111110000000000000011111111111110000000000000000011111111110000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111111111111000000000000000011111111111100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 832) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000010000000000000000000011100011100000000000000000001111111110000000000000001111111111110000000000011111111111111000000000000001110000111100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000111110000000000000001111111111111000000000000000111111111110000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 833) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001111111111111000000000000011111111111111100000000000011111111111111100000000000111111100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011111111111111000000000000001111111111111100000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 834) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000001111111111110000000000000000111111101111100000000000000111110000000110000000000000111100000000010000000000000011100000000000000000000000001111000000000000000000000000011110000000000000000000000000111111000000000000000000000001111111000000000000000000000011111110000000000000000000000111111000000000000000000001111110000000000000000000111111000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011111111000011000000000000000111111111111100000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 835) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000000000000000000000111111110000000000000000001111111111111100000000000001111100000111110000000000001111000000000000000000000000111000000000000000000000000011000000000000000000000000001110000000000000000000000000011110000000000000000000000000111111000000000000000000000000111111000000000000000000000000111100000000000000000000000011110000000000000000000000111110000000000000000000001111100000000000000000000011111100000000000000000000011110000000000000000000000011110000000000000000000000001111111111111100000000000000011111101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 836) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000001111111111100000000000000001111111111100000000000000001111110000000000000000000000111100000000000000000000000001111110000000000000000000000011111110000000000000000000000011111110000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000011100000000000001110000000001110000000000001111000000111111000000000000111111111111110000000000000001111111111100000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 837) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000110000000000000001111000000011100000000000000111100000001110000000000000111110000000111000000000000011111000111111100000000000001111111111111110000000000000111111111111111000000000000001111100001111100000000000000000000000011111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 838) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111110000000000000000111111111111000000000000000011110000000000000000000000000111110000000000000000000000001111110000000000000000000000001111111100000000000000000000011111111000000000000000000000001111110000000000000000000001111110000000000000000000001111100000000000000000000001111100000000000000000000000111111111111110000000000000111111111111111000000000000001110000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 839) begin
            pixels = 784'b0000000000000000000000000000000000000011100000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011111000000000000000000000001111100000000000000000000001111100000000011000000000000111110000010011110000000000011111011111111111100000000001111111111111111110000000000011111111111111111100000000000111110000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 840) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000011111111111000000000000000011111111111110000000000000011111000111111000000000000011111000000000000000000000001111100000000000000000000000111110000000000000000000000001111111110000000000000000000111111111110000000000000000001111111111000000000000000000001111111100000000000000000000011111100000000000000000000011111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000110000000000000000111111111111110000000000000001111111111111000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 841) begin
            pixels = 784'b0000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000000111110000000000000000000000011111000000000000000000000001111100000000000000000000000111100000000010000000000000111110000000001100000000000011111001111001111000000000001111111111111111100000000000111111111111111111000000000001111110000011111100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 842) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000001111111110000000000000000001111111111100000000000000000111111111110000000000000000011100000001000000000000000001110000000000000000000000000011100000000000000000000000001111100000000000000000000000011111100000000000000000000000011111100000000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000000011100000001100000000000000001111111111111000000000000000001111111111100000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 843) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000001000000000000001110000000001110000000000001111111111111111000000000000111111111111111100000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 844) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000011111111111111100000000000011111111111111110000000000011111110000000000000000000001111000000000000000000000000111000000000000000000000000001110000000000000000000000000011110000000000000000000000000111111111000000000000000000000111111100000000000000000000000111110000000000000000000000011111000000000000000000000011110000000000000000000000011111000000000000000000000011110000000000000000000000001111000000000110000000000000111100000000111100000000000001111111111111110000000000000001111111111100000000000000000001111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 845) begin
            pixels = 784'b0000000000000000000000000000000000000110000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000001100000000000011110000000001110000000000001111000000000111100000000000111100000111111110000000000111111111111111111000000000011111111111111111100000000001111111111111011110000000000011111000000000111000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 846) begin
            pixels = 784'b0000000000000000000000000000000000000011000000000000000000000000001110000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000011100000000000001111111100001110000000000000111111111100111100000000000011111111111111111000000000000111100001111111100000000000000000000011111110000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 847) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000111111100000000000000000001111111111100000000000000001111111111111110000000000001111111111111111100000000000111111100000111111000000000001111100000000111100000000000011110000000000110000000000001111100000000000000000000000011111100000000000000000000000011111000000000000000000000011111110000000000000000000011111111000000000000000000001111111100000000000000000000111111000000000000000000000011111000000000000000000000001111111111111000000000000000111111111111110000000000000000111111111111000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 848) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001111111001111110000000000001111111111111111100000000001111000111111110000000000000111100000000000000000000000001110000000000000000000000000111100000000000000000000000001111000000000000000000000000011111110000000000000000000000111111110000000000000000000000111111000000000000000000000111111100000000000000000000111111000000000000000000000111110000000000000000000000011110000000000000000000000001110000000000000000000000000111110000000110000000000000001111111111111000000000000000001111111111110000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 849) begin
            pixels = 784'b0000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000001000000000000000011100000001110000000000000001110000000011000000000000000111011111011100000000000000111111111111110000000000000111111111111111000000000000111111000011111100000000000011110000000011110000000000001100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 850) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000110000000000000001110000000011100000000000001111000000001100000000000000011100000000110000000000000011111111111111000000000000011111111111111100000000000001111111111111111000000000000111111100001111100000000000000100000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 851) begin
            pixels = 784'b0000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000001100000000000000011110000001111000000000000001110000000011100000000000000111000000001110000000000000111100011111111000000000000011111111111111100000000000001111111111111111000000000000011111000011111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 852) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000011111111111110000000000000001111111111111100000000000000111111111111111100000000000011000000000000010000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000001111000000000000000000000000011110000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001111000110000000000000000000011111111000000000000000000001111111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 853) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000111111111100000000000000001111111111111100000000000001111111111001100000000000000111110000000000000000000000011110000000000000000000000000111110000000000000000000000001111110000000000000000000000011111111000000000000000000000011111100000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000010000000000111110000000011111100000000011111111111111111100000000000111111111111111100000000000001111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 854) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000001111111111000000000000000001111111111100000000000000001111111111111000000000000000111111000011100000000000000011110000001110000000000000001111100000100000000000000000011111111000000000000000000000011111110000000000000000000000111111000000000000000000000011111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000000011100000000000100000000000001111111111001111000000000000011111111111111110000000000000111111111111110000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 855) begin
            pixels = 784'b0000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011110000000010000000000000011111000000011100000000000001111000000001110000000000000111100000000111000000000000011111111111111100000000000001111111111111111000000000000111111111111111100000000000011111101111111111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 856) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000011000000000000001111000000011100000000000000111111100001111000000000000011111111111111100000000000001111111111111110000000000000111111111111111100000000000000000000000111110000000000000000000000000111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 857) begin
            pixels = 784'b0000000000000000000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011111000001100000000000000001111100000110000000000000000111100000011100000000000000111110000001111000000000000011111000000111100000000000001111111111111110000000000001111111111111111000000000000111111110001111100000000000001111000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 858) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000111110000011100000000000000011110000001110000000000000001111000000111100000000000001111111110011110000000000000111111111111111000000000000011111111111111100000000000000111000001111110000000000000000000000001111000000000000000000000000011100000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 859) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111110000000000000000011111111111100000000000000011111111111110000000000000011111111000000000000000000000111110000000000000000000000001111000000000000000000000000011111000000000000000000000000111111000000000000000000000001111100000000000000000000001111111000000000000000000000111110000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000011110000000111100000000000000111100011111110000000000000001111111111111000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 860) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000001111111111000000000000000011111111111110000000000000011111111111111100000000000011111100000000110000000000001111000000000000000000000000011100000000000000000000000001111111110000000000000000000011111111110000000000000000000011111111000000000000000000000011111100000000000000000000011111110000000000000000000011111100000000000000000000011111000000000000000000000001111000000000000000000000000111100000000000000000000000001111000000000000000000000000001111111100000000000000000000011111111000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 861) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000001111111000000000000000000011111111100000000000000000011110000110000000000000000011110000000000000000000000011100000000000000000000000001110000000000000000000000001110000011100000000000000000111000111110000000000000000001111111110000000000000000000111111110000000000000000000001111100000000000000000000000111100000000000000000000000111100001100000000000000000111100011111000000000000000011100111111000000000000000001111111111000000000000000001111111110000000000000000000111111000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 862) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000110000000000000000011100000111100000000000000011100000011100000000000000011100000011100000000000000011111100111100000000000000011111111111100000000000000011111101111110000000000000011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 863) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000011111111111110000000000000111111110011111000000000000111110000000011000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000011100000011100000000000000001111111111110000000000000000011111111110000000000000000001111111000000000000000000001111110000011000000000000001111100000111100000000000000111000011111110000000000000011111111111100000000000000001111111110000000000000000000011111100000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 864) begin
            pixels = 784'b0000000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000001000000000000000111100000011110000000000000111100000011111000000000000111100000011111000000000000111111100111111000000000000111111111111111000000000000111110111111111000000000000001000000111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 865) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000001111111000000000000000000111111111000000000000000001111111110000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000011111111000000000000000000001111111100000000000000000001111110000000000000000000001111000000000000000000000001111101111110000000000000000111111111111000000000000000001111111111000000000000000000111111110000000000000000000111111100000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 866) begin
            pixels = 784'b0000000000000000000000000000000000000000000000011100000000000000000000000001111000000000000000000000011111000000000000000000000001111000000000000000000000011111000000000000000000000011111000000000000000000000011110000000000000000000000001111000000000000000000000011110000000000000000000000001111000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000011100000000000001111000000011110000000000001111000000111110000000000001111111111111110000000000001111111111111110000000000000011100000011110000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 867) begin
            pixels = 784'b0000000000000000000000000000000000000000000000111000000000000000000000001111100000000000000000000001111110000000000000000000000111110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000001110000000000000000000000001111000000000000000000000001110000000110000000000000001111000000111000000000000001111000000111100000000000001111000000111110000000000000111100000111110000000000001111000001111110000000000000111111111111111000000000000111111111111110000000000000011111111101111000000000000001111000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 868) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000111111111100000000000000001111111111110000000000000011111100001111000000000000011111000011111000000000000011110000000011000000000000001110000000000000000000000001110000110000000000000000000111111111000000000000000000011111111100000000000000000000111111000000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000011110000011110000000000000001110000111111000000000000000111011111111000000000000000011111111100000000000000000000111111100000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 869) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000111111111110000000000000001111111011111000000000000001111000001111000000000000011111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000001100000100000000000000000000111111111000000000000000000011111111100000000000000000011111110000000000000000000011111000000000000000000000011110000000000000000000000001110000011100000000000000001110000011110000000000000000111011111110000000000000000011111111110000000000000000000111111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 870) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000111111111110000000000000001111100000011100000000000001110000000001110000000000001110000001111111000000000000110000000001111000000000000011100000000000000000000000001111111110000000000000000000111111110000000000000000000011111100000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000011100001111000000000000000001111111111100000000000000000011111111000000000000000000000111110000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 871) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000111111111110000000000000001111110111111100000000000001111000000011100000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011110011000000000000000000001111111110000000000000000000011111111000000000000000000011111110000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000111000111110000000000000000011111111111000000000000000000111111110000000000000000000011111000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 872) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111110000000000000000011111111111000000000000000011110000111100000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100001111000000000000000001111111111100000000000000000011111111000000000000000000000111110000000000000000000000011110000000000000000000000001110001111000000000000000001110001111100000000000000000111111111000000000000000000011111111000000000000000000001111110000000000000000000000011100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 873) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001111111111110000000000000011111110011111000000000000011111000001111000000000000011110000000011000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000011000111100000000000000000001111111111000000000000000000011111111000000000000000000001111100000000000000000000001111000000000000000000000001110000000100000000000000001111000011111000000000000001111000111111100000000000000111111111111000000000000000011111111100000000000000000000111111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 874) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000001111111111111100000000000011111100000111100000000000011110000001111100000000000001110000000000000000000000001111000000000000000000000000111000011100000000000000000011100111110000000000000000001111111111000000000000000000011111111000000000000000000011111000000000000000000000011110000000000000000000000011110000011100000000000000001110000111110000000000000000111111111111000000000000000011111111100000000000000000000111111100000000000000000000001111000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 875) begin
            pixels = 784'b0000000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000011000000000000001111000000011100000000000001111000000011110000000000000111100000111110000000000000111111111111110000000000000011111111111111000000000000001111000001111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 876) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000001110000000000000000111000001111000000000000000111000001111100000000000000111000001111000000000000000111110001111100000000000000011111111111100000000000000011111111111100000000000000011111111111100000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 877) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111100000011000000000000000111100000011100000000000000111100000111110000000000000011111111111110000000000000011111111111110000000000000000111111011110000000000000000000000001110000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 878) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111110000000000000000111111111111100000000000000111100000111100000000000000111100000000110000000000000111100000000000000000000000001110000000000000000000000001111000000000000000000000000011111100011000000000000000000111111111110000000000000000001111111110000000000000000000111110000000000000000000000111100000000000000000000000011110000000000000000000000001100000011100000000000000000111111111110000000000000000011111111110000000000000000001111111110000000000000000000111111000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 879) begin
            pixels = 784'b0000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000011100000000000000111100000001110000000000000111100000001110000000000000011111000001111000000000000011111111111110000000000000001111111111111000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 880) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000110000000111110000000000000011101111111111000000000000001111111111101100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 881) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000111111000000000000000000001111101110000000000000000000111000001000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000000011000000000000000000000000001110000000000000000000000000011111100000000000000000000000111110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000000110001110000000000000000000011111110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 882) begin
            pixels = 784'b0000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000111011100000000000000111111111111111100000000000011111111111111110000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 883) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000111100000000000000000000000011000000000000000000000000011000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000011100000000000000000000000000111100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011111111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 884) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000001000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111111111111111100000000000011111111111111111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 885) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001111111111110000000000000000111111111111000000000000000000011111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 886) begin
            pixels = 784'b0000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000111000000000000000000111111111111110000000000000011111111111111000000000000000000010111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 887) begin
            pixels = 784'b0000000000111000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001111111111111111100000000001111111111111111110000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 888) begin
            pixels = 784'b0000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000001111111111110000000000000000111111111111111100000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 889) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111100000000000000000000111111111000000000000000000111100001100000000000000000111000001100000000000000000011000000000000000000000000001100000000000000000000000000100000000000000000000000000111000000000000000000000000001110000000000000000000000000011111100000000000000000000000111110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011110000110000000000000000000111111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 890) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000111111100000000000000000000111000011000000000000000000011000000100000000000000000001000000010000000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000001100000000000000000000000000110000000000000000000000000001100000000000000000000000000111000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000001000000000000000000000000000110000001000000000000000000001111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 891) begin
            pixels = 784'b0000000000000000000000000000000000000000010000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100011111111100000000000000111111111111110000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 892) begin
            pixels = 784'b0000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001111111111111111100000000000011111111111111111000000000000110111101000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 893) begin
            pixels = 784'b0000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000111111111111110000000000000011111111111111000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 894) begin
            pixels = 784'b0000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111011111111111000000000000001111111111111110000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 895) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000001111111000000000000000000011111111100000000000000000001111000010000000000000000001111000001100000000000000000111000000110000000000000000111000000010000000000000000011000000000000000000000000001100000000000000000000000000011000000000000000000000000001111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000001100000000000000000000000000111000011000000000000000000001111111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 896) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000111000000000000000001111111111111000000000000000011111111111110000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 897) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111100000000000000000111111000111000000000000000011110000000110000000000000011100000000001000000000000001100000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000000000000000000100000000000000000000000000001000000000000000000000000000110000000000000000000000000001110000000000000000000000000011000000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000011000100000000000000000000001111111000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 898) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111111000000000000000000011111111110000000000000000011110000011000000000000000001110000001100000000000000000110000000100000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000011000000000000000000000000001111000000000000000000000000011100000000000000000000000000110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000001100000000000000000000000000111100000000000000000000000001111111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 899) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111111000000000000000000011111111100000000000000000011111000011000000000000000011110000000100000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000000111110000000000000000000000001111100000000000000000000000011110000000000000000000000011111000000000000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001111000100000000000000000000011111110000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 900) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001111111000000000000000000001111111111000000000000000001111111111110000000000000000111000001111000000000000000111000000001100000000000000011000000000000000000000000001110000000000000000000000000011000000000000000000000000001111000000000000000000000000001111111000000000000000000000011111110000000000000000000000111111000000000000000000000111111000000000000000000000011110000000000000000000000001110000000000010000000000000111100000000111000000000000001111111111111100000000000000001111111111000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 901) begin
            pixels = 784'b0000000000001000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000001100000000000001111000000000110000000000001111000000000111000000000000111100000000111110000000000011111101100111110000000000001111111111111110000000000000011111111111111000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 902) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111100000000000000000011111111110000000000000000011111000000000000000000000011110000000000000000000000000110000000000000000000000000011110000000000000000000000000011110000000000000000000000000111111100000000000000000000000011111000000000000000000000001111100000000000000000000001111100000000000000000000001111000000000000000000000000011000000000111000000000000000111111111111000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 903) begin
            pixels = 784'b0000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000100000000000000111100000000010000000000000011110000000001000000000000011110000000001111000000000001111111111111111100000000000111111111111111100000000000001111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 904) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000011111111100000000000000000011111111110000000000000000111111000000000000000000000111110000000000000000000000011110000000000000000000000001111100000000000000000000000011111110111110000000000000000111111111111000000000000000000111111111000000000000000000000111111000000000000000000000011110000000000000000000000001110000000000000000000000000110000000000100000000000000011100000000111000000000000011111100000111000000000000000111111111111100000000000000001111111111100000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 905) begin
            pixels = 784'b0000000000000000000000000000000000000001110000000000000000000000000111100000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000110000000000001111000000000111000000000000111000000000011100000000000011100000000011110000000000011111111111111111000000000001111111111111111100000000000111111111111111100000000000001110011111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 906) begin
            pixels = 784'b0000000000000000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000110000000000000011100000000111100000000000001110000000011110000000000000111000000001111000000000000011100000000111100000000000001110000000011110000000000001111111111111111000000000000011111111111111100000000000000001111011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 907) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000001111111111111110000000000001111111111111111000000000001111111100000011000000000000111100000000000000000000000011100000000000000000000000001111110000000000000000000000011111111100000000000000000000011111111000000000000000000011111111100000000000000000111111111100000000000000000111111100000000000000000000011110000000000000000000000011110000000000000000000000001110000000011000000000000000111100000001110000000000000011111000001111000000000000000111111111111100000000000000001111111111100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 908) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000100000000000000000011100000110000000000000000011110000111000000000000000001111001111000000000000000000111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 909) begin
            pixels = 784'b0000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000001100000000000001110000010111110000000000000111111111111111000000000000001111111111111100000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 910) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000111111111000000000000000001111111101100000000000000001111100000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000000111100000000000000000000000001111111100000000000000000000001111111000000000000000000000111111100000000000000000000111111100000000000000000000111100000000000000000000001111000000000000000000000000110000000001000000000000000011000000000100000000000000001100000000110000000000000000111110011111000000000000000001111111111000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 911) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000011111111111000000000000000111111111111100000000000000111111111111110000000000000111100000000100000000000000011100000000000000000000000011110000000000000000000000000111110000000000000000000000001111111000000000000000000000011111111100000000000000000000011111110000000000000000000001111110000000000000000000001111100000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100001110000000000000000000111111111000000000000000000011111111000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 912) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000011111111000000000000000000111110000000000000000000000111100000000000000000000000011000000000000000000000000011100000000000000000000000000111000000000000000000000000001110000000000000000000000000111100000000000000000000000001111100000000000000000000000001111000000000000000000000000111100000000000000000000001111100000000000000000000001111100000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011111100100000000000000000000111111111000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 913) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000011111111000000000000000000111111111110000000000000001111111100011000000000000001111100000000000000000000001111000000000000000000000001110000000000000000000000000011100000000000000000000000001110000000000000000000000000011111111000000000000000000000111111110000000000000000000001111111000000000000000000000011111000000000000000000000011111000000000000000000000011110000000000000000000000001111000000000000000000000001111000011110000000000000000111111111111000000000000000001111111111000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 914) begin
            pixels = 784'b0000000000000000000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000001100000000000000000011000000110000000000000000001100000011000000000000000000111100001100000000000000000001111110110000000000000000000001111111000000000000000000000000111100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 915) begin
            pixels = 784'b0000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000001000000000000000000110000000100000000000000000011000000110000000000000000001111111111000000000000000000111111111000000000000000000000001011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 916) begin
            pixels = 784'b0000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000110000000000000011000000000011000000000000001111000000001100000000000000111111111001110000000000000000011111111111000000000000000000000011111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 917) begin
            pixels = 784'b0000000000000000000000000000000000000001111000000000000000000000000011110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000001000000000000001110000000001110000000000000110000000001111000000000000111000000000111000000000000011100000000111000000000000001100000000011100000000000000111110000111110000000000000001111111111110000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 918) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111100000000000000000111111111110000000000000001111110000000000000000000001111100000000000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000001111000000000000000000000000011111100000000000000000000000111110000000000000000000000111111000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001110000000011100000000000000011111111111100000000000000000111111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 919) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000110000000000000000000110000011000000000000000000111000001110000000000000000011100000111000000000000000000110000001100000000000000000011000000110000000000000000001111101111100000000000000000011111111110000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 920) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000111111111110000000000000001111111111111100000000000001111111111111100000000000000111111000000010000000000000011110000000000000000000000001111100000000000000000000000011111111100000000000000000000111111110000000000000000000011111111000000000000000000111111111000000000000000000111111100000000000000000000111111000000000000000000000011110000000000000000000000001110000000000000000000000000111100000000000000000000000001111110110000000000000000000011111111100000000000000000001111111110000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 921) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000010000000001110000000000000001000000001111000000000000000000000000111000000000000000010000000111000000000000000001000000011100000000000000000100000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000110000000000000001110000000011000000000000000111000000011100000000000000011111111111110000000000100001111111111110000000000010000011111111110000000000001000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 922) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000001111111000000000000000000011111111110000000000000000011110000011000000000000000011110000001100000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000000110000000000000000000000000011100000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100010000000000000000000001100011100000000000000000000011111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 923) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111111000000000000000000111111111100000000000000001111111111110000000000000001111110000100000000000000001111100000000000000000000000111100000000000000000000000001111000000000000000000000000011111000000000000000000000001111100000000000000000000011111110000000000000000000011111110000000000000000000011111000000000000000000000011111000000000000000000000001110000000000000000000000001110000001000000000000000000011000001110000000000000000001111111111000000000000000000011111111000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 924) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011111111000000000000000000001111111111111100000000000000001111111111110000000000000000000000111111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 925) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000011111000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000011100001110000000000000000001111111111100000000000000000011111111110000000000000000000011111110000000000000000000001111100000000000000000000001111110000000000000000000000111111100000000000000000000011111111111100000000000000000111111111111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 926) begin
            pixels = 784'b0000000000000000000000000000000000000011100000000000000000000000001111000000000000000000000000111000000000000000000000000001110000000000000000000000001110000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000001111000000000000000000000000111100000000000000000000000011111110000000000000000000001111111111100000000000000000111111111111000000000000000000111111111110000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 927) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000011110000000000000000000000111111000000000000000000001111110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000000111100000000000000000000000011110000000000000000000000001111111100000000000000000000011111111000000000000000000000111111100000000000000000000011111110000000000000000000011111110000000000000000000011111000000000000000000000001111100000000000000000000000111111111110000000000000000001111111111100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 928) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111111000000000000000000000000011110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011111000000000000000000000001110000000000000000000000000111111100000000000000000000011111111110000000000000000000011111111110000000000000000000001111111100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 929) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000111111111000000000000000000111111111100000000000000001111111000110000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011111000000000000000000000001111111000000000000000000000011111111100000000000000000000111111110000000000000000000011111110000000000000000000011111100000000000000000000011111110000011000000000000000111111111111100000000000000001111111111110000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 930) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000011110000000000000000000000000111100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000001111100000000000000000000000111100000000000000000000000011110000000000000000000000011111000000000000000000000001111011000000000000000000001111111111100000000000000000111111111111100100000000000011111011111111110000000000000000000000111111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 931) begin
            pixels = 784'b0000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000000111100000001100000000000000111110000001110000000000000011110000001111000000000000011110000001111100000000000001111000001111110000000000000111100011111110000000000000011110111111111000000000000001111111111011000000000000000111111110000000000000000000011111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 932) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111000000000000000000001111111100000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000000111100000000000000000000000011111111000000000000000000000011111110000000000000000000001111110000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001111000000000000000000000000011110010000000000000000000000111111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 933) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011111000000000000000000000001111000000110000000000000000111100000111100000000000000011100000011100000000000000001110000011110000000000000000110000001110000000000000000011000000110000000000000000001111111111000000000000000000111111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 934) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111100000000000000000000011111110000000000000000000001110010000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111111110000000000000000000011111111000000000000000000001111111100000000000000000000111111100000000000000000000111110000000000000000000000111100000000000000000000000011100000100000000000000000001111100111000000000000000000111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 935) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000100000000000000011110000001111000000000000001110001111111100000000000000111111111111110000000000000011111111110111000000000000000111110000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 936) begin
            pixels = 784'b0000000000000001100000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000110000000000000001110000000111000000000000011110000001111100000000000001111000001111100000000000000111000001111100000000000001111111111111110000000000000111111111111110000000000000001111111111110000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 937) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000111111111100000000000000000111111111110000000000000000111110000011000000000000000011110000011100000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000001111101111110000000000000000111111111111000000000000000001111111111000000000000000001111111000000000000000000011111111000000000000000000001111110000000000000000000000111110000000000000000000000011111100000000000000000000000111111110011000000000000000000111111111100000000000000000000011111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 938) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000111111111000000000000000000111110011100000000000000000111100000010000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111100000000000000000000000001110000000000000000000000000111100000000000000000000000001111111110000000000000000000011111111000000000000000000011111111100000000000000000111110100000000000000000001111110000000000000000000000111100000000000000000000000011110000000000000000000000001111111111100000000000000000011111111110000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 939) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111100000000000000000000111111111000000000000000001111000001000000000000000001111000000100000000000000001110000000000000000000000000110000000000000000000000000011000001000000000000000000011100111100000000000000000001111111110000000000000000000111111100000000000000000000011111000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000000000000000000000001111000100000000000000000000011111111100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 940) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111111111000000000000000000011111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 941) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000001111111000000000000000000001111111100000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001111111111110000000000000000011111111110000000000000000001111111100000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000011110000001100000000000000001111111111110000000000000000011111111111100000000000000000001111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 942) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000001111000000000000000000000000011100000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000000111100000000000000000000000011110000000000000000000000111110000000000000000000000011110000001110000000000000011111111111111100000000000011111111111111110000000000001111111111111111000000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 943) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000001100000000000111110000000001110000000000011110000111111110000000000001111111111111111000000000000111111111111110000000000000011111111111100000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 944) begin
            pixels = 784'b0000000000000000000000000000000000000000001110000000000000000000000001111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000001111100000000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111110000000001000000000000011111111111111111100000000001111111111111111110000000000110000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 945) begin
            pixels = 784'b0000000000000000000000000000000000000000001100000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000110000000000000000001110000111000000000000000000111000111100000000000000000011110111110000000000000000001111111110000000000000000000111111110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 946) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111100000000000000000111111111100000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111111100000000000000000000001111111111000000000000000000011111111100000000000000000000011111110000000000000000000011111000000000000000000000011111000000000000000000000011111000010000000000000000001111110111000000000000000000111111111100000000000000000000111111110000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 947) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000001111111000000000000000000011111111000000000000000000011110000000000000000000000111110000000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111111011111000000000000000001111111111100000000000000000001111111100000000000000000000111110000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001111000000000000000000000000111111111100000000000000000001111111111000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 948) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000001111111111000000000000000011111111111100000000000000011111100000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000011111110000000000000000000000111111000000000000000000000111111000000000000000000000011111000000000000000000000011111000000000000000000000001111111000000000000000000000011111110000000000000000000000011111100000000000000000000000001111000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 949) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011110000000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000001111100000000000000000000001111100000000000000000000001111100000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011100000000000000000000000001111000000000000000000000000111111000000000000000000000011111111111110000000000000000111111111111100000000000000001111111111110000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 950) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000011111111111111000000000000111111111111111110000000000111110011111111111000000000111100000000000000000000000011100000000000000000000000000110000000000000000000000000011100000000000000000000000000111000000000000000000000000001111100000100000000000000000001111111111000000000000000000001111111000000000000000000000111100000000000000000000001111000000000000000000000011111000000000000000000000011111000000000000000000000011110000000000110000000000001110000000111111100000000000111111111111111110000000000000111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 951) begin
            pixels = 784'b0000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000111110000000000000000000000111111000000000000000000000011110000000000000000000000011111000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111100000000000000000000000011110001111111110000000000001111111111111111100000000000011111101001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 952) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000111111111110000000000000001111111111111100000000000000111111111111111000000000000111100000011111100000000000011100000000001000000000000011110000000000000000000000000111000000000000000000000000001110000000000000000000000000111100000000000000000000000001111111110000000000000000000011111111000000000000000000011111111100000000000000000111111111000000000000000011111100000000000000000000001111000000000000000000000001111000000000000000000000000111100001110000000000000000001111111100000000000000000000011111000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 953) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000111110000000000000000000000011100000000000000000000000011110000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000001110000000000001110000001111111000000000000111000111111111110000000000001111111111000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 954) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000001111111111000000000000000001111111111110000000000000001110000001111000000000000000111000000000000000000000000001110000000000000000000000000011100000000000000000000000000111000000000000000000000000001111100000000000000000000010011111000000000000000000001101111100000000000000001001111110000000000000000000111111000000000000000000000011110000000000000000000000111100000000000000000000000111100000000000110000000000011100000000011111100000000001110000000111101100000000000011101110010000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 955) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000111100000000000000000000000111100000000000000000000001111100000000000000000000000100000000000000000000000000011100000000000000000000000011100000000000000000000000111100000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000100001111111110000000001101111111111111111000000000000000001111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 956) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111011100000000000000000000111111100000000000000000000111101101111111110000000000110000000000001110000000000011000000000000000000000000000110000000000000000000000000011000000000000000000000000000110011000000000000000000000001111100000000000000000000000011100000000000000000000000001110000000000000000000000000100000000000000000000000001100000000000000000000000001100000010000000000000000011110011100011100000000000011110011000011110000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 957) begin
            pixels = 784'b0000000000000000000000000000000000000000000000001000000000000000000000001111000000000000000000000001111000000000000000000000011110000000000000000000000011111000000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000001111000000000011111111110000111000000000001111111000111111100000000000011000011111111000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 958) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000001111000000000000000000000001111000000000000000000000000100000000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000100000000000000011100001111111000000000000001111111110111100000000000000011100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 959) begin
            pixels = 784'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000110000000000000011100000111111000000000000000111111111100000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 960) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000001111000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000111100000000000000000000000011110000000000000000000000011100000000001100000000000001110000000011111000000000011110000000011111000000000001110000000011110000000000001111111110111110000000000001111111111111110000000000000111111000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 961) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000111000000000000000000000001111000000000000000000000001111000000000000000000000001111000000000000000000000011110000000000000000000000011110000000000000000000000111110000000000000000000000011110000000000000000000000111110000000000000000000000111100000000000000000000000111100000000000000000000000011100000000111000000000000011110000000111100000000000011110000001111100000000000001110000001111100000000000000011100001111100000000000000001111111111100000000000000000000011111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 962) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000001111111111110000000000000011111000000011100000000000001110000000000010000000000000011000000000000000000000000000110000000000000000000000000001100000000000000000000000000011000000000000000000000000011110000000000000000000000011100000000000000000000000111100000000000000000000001111100000000000000000000001111000000000000000000000001111000001110000000000000001111000111111000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 963) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000001111110111100000000000000011110000000000000000000000011100000000000000000000000001100000000000000000000000000010000000000000000000000000000100000000000000000000000000001110000000000000000000000011001000000000000000000001110000000000000000000000011100000000000000000000000111100000000000000000000000011110001110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 964) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000011111111111111100000000000011111111111111100000000000011100000000000000000000000000110000000000000000000000000011000000000000000000000000000110000000000000000000000000001100000000000000000000000000011100000000000000000000000011110000000000000000000000111100000000000000000000011110000000000000000000000011100000000000000000000000001100000001000000000000000000011111111110000000000000000000111011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 965) begin
            pixels = 784'b0000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000111110000000000000000000000111100000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000111000000000001110000000000111100000000001110000000000111100000000001110000000000111100000000000111000000000111100000000000111000111111111100000000000011111111111111100000000000000110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 966) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000001111111111111000000000000000011111111111110000000000000001110000000001000000000000000011000000000000000000000000001110000000000000000000000000011100000000000000000000000000011100000000000000000000000011110000000000000000000000111000001100000000000000001110000000000000000000000011100000000000000000000000011000000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000110000000000000000000111111111100000000000000000011111111111000000000000000000010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 967) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000001111110000000000000000000011111111100000000000000000011110000011100000000000000001100000000110000000000000000110000000000000000000000000011000000000000000000000000000000000000000000000000000000011001000000000000000000000000111111000000000000000000000111111100000000000000000001111000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001110000001100000000000000000110000001110000000000000000110001111111000000000000000001111111110000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 968) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111100000000000000000000111111000000000000000000000011000000110000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000011110000000000000000000000000111100000000000000000000000011100000000000000000000000011000000000000000000000000111000000000000000000000000111000000000000000000000000110000000010000000000000000110000000011100000000000000011000000111111000000000000001100001111110000000000000000001111110000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 969) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111000000000000000000000000111000000000010000000000000111100000000011100000000000011100000000011110000000000011100000000011110000000000001110000000011110000000000001110000000011111000000000001110000000011111000000000000111100011111111000000000000011111111111111100000000000000111111100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 970) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000001001000000000000000000000000101000000000000000000000000001100000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000001100000000000001110000000011110000000000000111000000011000000000000000111000000000000000000000000011100000000011100000000000001111111111011100000000000000111111001111110000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 971) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101000000000000000000001111110011000000000000000111111111111100000000000001111110000111100000000000011111100000000000000000000001111000000000000000000000000011100000000000000000000000000111100000000000000000000000000011100000000000000000000000000011110000000000000000000000000111100000000000000000000000111110000000000000000000011110000000000000000000000011110000000000000000000000111100000000000000000000000111100000000010000000000000111000000000111100000000000011100000000110100000000000000111100011000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 972) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000001111111111111110000000000001111101000011111100000000001111100000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000001110000111000000000000000000111101111110000000000000000001111111111000000000000000000011111111100000000000000000001111111100000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000001110000000000000001110000001110000000000000000011100111110000000000000000001111111111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 973) begin
            pixels = 784'b0000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100001100000000000000000011100000110000000000000000001100000110000000000000000011100000111000000000000000001110000011000000000000000001110000011100000000000000001111111111100000000000000001111111111110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 974) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111111111000000000000001111000000111110000000000001110000000000111100000000000111000000000001110000000000111000000000000000000000000011100000000000000000000000001110000110000000000000000000011001111100000000000000000001111111110000000000000000000111110011000000000000000000011111111000000000000000000001111111000000000000000000000110010000010000000000000000111000000011000000000000000011100000001100000000000000001110000011110000000000000000011110111110000000000000000000111111110000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 975) begin
            pixels = 784'b0000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000011000000000000000001110000011100000000000000001110000011100000000000000011111000001100000000000000011111111001110000000000000001111111111110000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 976) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111110000000000000001111110000001000000000000011111000000000100000000000011110000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011100011111000000000000000000111111111100000000000000000011111101110000000000000000001111111110000000000000000000111001110000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011100001100000000000000000001111111110000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 977) begin
            pixels = 784'b0000000000000000000000000000000000000000000000001100000000000000000000000011110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000100000000000000000011100000110000000000000000011000000011000000000000000111000000111000000000000000111000000111000000000000000111100000011100000000000001111000000011100000000000001111111110111100000000000000111111111111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 978) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000010000000000000000001110000011100000000000000001110000011100000000000000001110000001110000000000000000111000001110000000000000000111000000111000000000000000011111111111000000000000000001111111111000000000000000000011111111100000000000000000000000001110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 979) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000111111111000000000000000011111110001110000000000000011110000000011100000000000011100000000000110000000000011100000000000011000000000001100001111000011100000000001110000001111111100000000000111000011000000000000000000011100111110000000000000000000111111111000000000000000000011111111100000000000000000011111111100000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000000111000000000000000000000000001111000000000000000000000000011111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 980) begin
            pixels = 784'b0000000000000000000000000000000000000000000000001000000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000110000000000000000001100000111000000000000000001100000011000000000000000001110000011000000000000000001111111011000000000000000011111111111100000000000000001111000001100000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 981) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000011000000000000000000110000001100000000000000000110000001110000000000000000111000001111000000000000000011000001111100000000000000011000000111100000000000000011111111111100000000000000001111110111110000000000000000100000001110000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 982) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000001000001111111111100000000001100001111101111111100000000110001110000000111110000000011001111000000000110000000001101111000000000000000000000110111000000000000000000000011011100000000000000000000001101110001100000000000000000110111011111000000000000000011001111111100000000000000001000111101110000000000000000000111111110000000000000000000011111110000000000000000000011100000000000000000000000101110000010000000000000000011111000011000000000000000001101111111100000000000000000000111111100000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 983) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001111110000000000000000000011110001100000000000000000011100000011000000000000000011100000111100000000000000001100000001100000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000001100000011000000000000000000110000111100000000000000000011111111110000000000000000000111111111000000000000000000001111100000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000011000011000000000000000000001111111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 984) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111100000000000000000000111000010000000000000000000110000001000000000000000000110000001100000000000000000010000001100000000000000000011000001100000000000000000001000000000000000000000000001100000100000000000000000000110001111000000000000000000011001111000000000000000000001101111000000000000000000000011110000000000000000000000001100000000000000000000000000100000000000000000000000000110000000000000000000000000110001000000000000000000000011001100000000000000000000000111110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 985) begin
            pixels = 784'b0000000000000000000100000000000000000000000000110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000110000011100000000000000000110000011100000000000000000111000001110000000000000000111000001110000000000000000011111111110000000000000000001111001111000000000000000000000000111000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 986) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000001110000001000000000000000001110000001110000000000000000110000000111000000000000000111000000111000000000000000111000000111000000000000000011000000111000000000000000011000000111000000000000000001111111111000000000000000001111111111100000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 987) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000001110000000000000000000000000111000000100000000000000001111000001110000000000000001111000001111000000000000000111000000111000000000000000111100000111000000000000000111111111111000000000000000111111111111100000000000000011100000111100000000000000000000000011100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 988) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000111000000000000000000000000111000000100000000000000000111000000110000000000000000111000000111000000000000000111000000111000000000000000111000000111000000000000001111000001111000000000000001111100011111100000000000000011111111111100000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 989) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111111100000000000000011110000000110000000000000011110000000001000000000000001110000000001100000000000001110000000000100000000000000111000000000000000000000000011100000000000000000000000000110000110000000000000000000011111111000000000000000000000111111100000000000000000000111111110000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001111100000000000000000000000001111111000000000000000000000000111100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 990) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000011000000000000000111000000011100000000000000011000000011100000000000000011110000111100000000000000011111111111000000000000000000000011111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 991) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111111000000000000000000111110000110000000000000000111100000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000010000000000000000000011000111100000000000000000001111111100000000000000000000011111000000000000000000000000111000000000000000000000000011000000000000000000000000011100001100000000000000000001110001110000000000000000000011111110000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 992) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000001111111110000000000000000001111111111100000000000000011110000000011000000000000001110000000001100000000000001110000000000000000000000000110000000000000000000000000111000110000000000000000000011101111100000000000000000000111111100000000000000000000011110110000000000000000000001111110000000000000000000000111111000000000000000000000011110000000000000000000000011000000100000000000000000001100000110000000000000000000110001110000000000000000000011101110000000000000000000000111110000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 993) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000111111111100000000000000000111111111111000000000000000111110011111100000000000000011100000111110000000000000011100000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000001110000000000000000000000000011111100000000000000000000000111110000000000000000000000111110000000000000000000000111110000000000000000000000111100011100000000000000000111100011110000000000000000011111111110000000000000000001111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 994) begin
            pixels = 784'b0000000000000000000000000000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000110000000000000000001111111111110000000000000000011111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 995) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000111111100000000000000000001111111111000000000000000001111001111100000000000000001110000011110000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000001000000000000000000000000000110000010000000000000000000011100111000000000000000000000111111100000000000000000000001111110000000000000000000001111000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000011000111000000000000000000000111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 996) begin
            pixels = 784'b0000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000001000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011100111100000000000000000000111111111000000000000000000011111111000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 997) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111100000000000000001111111111111000000000000001111111001111110000000000001111100000001111000000000001111000000000011100000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000111000011100000000000000000001111111111000000000000000000011111111000000000000000000000111111000000000000000000000111110000000000000000000000011110000000000000000000000001110000000000000000000000000111000011100000000000000000011111111111000000000000000000111111111000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 998) begin
            pixels = 784'b0000000000000000000000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001111111111000000000000000000111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 999) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000011111111000000000000000000011111111110000000000000000001100000111100000000000000001100000000110000000000000001100000000001000000000000000110000000000000000000000000010000000000000000000000000001000000000000000000000000000100000100000000000000000000010001111000000000000000000001101111100000000000000000000111111110000000000000000000001111110000000000000000000000111100000000000000000000000110001100000000000000000000011001110000000000000000000001111111000000000000000000001111110000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1000) begin
            pixels = 784'b0000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000001000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011100101100000000000000000000111111111000000000000000000011111111100000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1001) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000001111111100000000000000000011111111110000000000000000011111111111000000000000000011000111111100000000000000011000000011100000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000111000000000000000000001111111000000000000000000000011111000000000000000000000001110000000000000000000000000110000100000000000000000000010000110000000000000000000011111111000000000000000000001111111000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1002) begin
            pixels = 784'b0000000000000000100000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000110000000000000011111111111111000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1003) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000000100000000000000000000000000110000000000000000000000000010000000000000000000000000010000000000000000000000000011000000000000000000000000001000000000000000000000000001100000000000000000000000000100000000000000000000000000110000000000000000000000000010000000000000000000000000001000000000000000000000000001000000000000000000000000000100000000000000000000000000100000000000000000000000000010000000000000000000000000010000000000000000000000000011000000000000000000000000001111111111110000000000000000111110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1004) begin
            pixels = 784'b0000000000000000000000000000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000011000000000000000110000001111100000000000000111000011111110000000000000011111111111100000000000000001111111110000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1005) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001111111111100000000000000001111100111111000000000000001110000000011110000000000000110000000000011000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000000100000000000000000000000000011101111000000000000000000000111111110000000000000000000011111111000000000000000000011110000000000000000000000001100000000000000000000000001110000000000000000000000000111001111100000000000000000001111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1006) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000001100000000000000000011001111111000000000000000011111111111000000000000000001111111100000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1007) begin
            pixels = 784'b0000000000000000000000000000000000000000000000100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000001111000000000000000011011111111100000000000000001111111110000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1008) begin
            pixels = 784'b0000000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000111110000000000000110000111111111000000000000111111111111111000000000000011111111100000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1009) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111110000000000000001111111111111000000000000001111100111111000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001110000000000000000000000000011100000000000000000000000000111111111100000000000000000001111111110000000000000000000001111110000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000001110000010000000000000000000011111111000000000000000000000111111100000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1010) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000111111100000000000000000000011111111000000000000000000011000111100000000000000000011000000110000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000011000000000000000000000000001111010000000000000000000000001111100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110011000000000000000000000111111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1011) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000111111000000000000000000000111111100000000000000000000111011110000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000100000000000000000000000000010000000000000000000000000001100000000000000000000000000111100100000000000000000000001111111000000000000000000000011111100000000000000000000000111100000000000000000000000011100000000000000000000000001100100000000000000000000001100111000000000000000000000111111100000000000000000000011111100000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1012) begin
            pixels = 784'b0000000000000000000000000000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000010000000000000000000000000011000000000000000000000000001100000011000000000000000001100000111110000000000000000110001111100000000000000000111011110000000000000000000011111100000000000000000000001111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1013) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000011111110000000000000000000011100000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000001000000000000000000000000000110000000000000000000000000011111100000000000000000000000111110000000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000001110010000000000000000000000011111100000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1014) begin
            pixels = 784'b0000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000001100000000000000000000000001110000111100000000000000000110111111110000000000000000011111111100000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1015) begin
            pixels = 784'b0000000000000000000000000000000000000000000000100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000001110000000111000000000000000110000011111100000000000000111011111111000000000000000011111111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1016) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000011110000000000000000000000011110000000100000000000000001110001111111110000000000000111001111111111000000000000011111111100111100000000000000111100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1017) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100011000000000000000000000111111100000000000000000000011111110000000000000000000011111110000000000000000000111100000000000000000000000111100000000000000000000000111100000000000000000000000111000000000000000000000000011100000000000000000000000001111111111100000000000000000001111111110000000000000000000000011100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1018) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000001100000000000000111000000111111000000000000011100000111111000000000000001100011111111000000000000000111111110110000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1019) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111111000000000000000000011110001110000000000000000011100000111000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000001100000000000000000000000000110000000000000000000000000011001110000000000000000000001111111000000000000000000001111110000000000000000000011110000000000000000000000011110000000000000000000000001110000111000000000000000001111111111100000000000000000011111111110000000000000000000000001110000000000000000000000011100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1020) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000011100000000001110000000000001110000000001111100000000001111000000001111100000000000111000000011111000000000000001100000011110000000000000000111110011100000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1021) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011100000011000000000000000011100000011100000000000000001110000011110000000000000001110000111100000000000000000111000011100000000000000000111111111100000000000000000011111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1022) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000011111111110000000000000000111110111110000000000000000110000000000000000000000000011000000000000000000000000011000010000000000000000000001100011100000000000000000000111111110000000000000000000011111100000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000011100000011000000000000000011100111111100000000000000011111111111100000000000000001110001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1023) begin
            pixels = 784'b0000000000000000000000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000011100000000000011100000000011100000000000001100000000111100000000000001110000000111100000000000000111110000111000000000000000111111111111000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1024) begin
            pixels = 784'b0000000000000000000000000000000000000000000011000000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000001100000000000000000011001111111000000000000000001111111110000000000000000000111111000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1025) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000001111111111100000000000000001111111111111000000000000001111100000011110000000000001111000000000110000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000011110000000000000000000000000111111110000000000000000000001111111100000000000000000000011111100000000000000000000111111000000000000000000001111110000000000000000000001111110000000000000000000001111000000011000000000000001111111111111000000000000001111111111111000000000000000111111111100000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1026) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000001111111110000000000000000001110000011100000000000000001100000001110000000000000000110000000111000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011000011100000000000000000001111111110000000000000000000011111110000000000000000000000111000000000000000000000000110000000000000000000000000111000001110000000000000000111000001111000000000000000111000011111000000000000000011001111111000000000000000011111111111000000000000000011111000010000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1027) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000101111111000000000000000001110000001000000000000000001110000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001111101110000000000000000000011111111000000000000000000000011111100000000000000000000001111000000000000000000000001111000011000000000000000001010000111100000000000000011100000111110000000000000011110000111100000000000000001100001111000000000000000011110011111000000000000000001111111111000000000000000001111111111000000000000000000011111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1028) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011100000001100000000000000011100000001110000000000000001110000001110000000000000001111000011110000000000000000000111111110000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1029) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000011100111111000000000000000001111111111100000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1030) begin
            pixels = 784'b0000000000000000000000000000000000000000000001000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000000000000000000000110000000000000000000000000110000000000000000000000000110000000000000000000000000110000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000100000000000000011100000011111000000000000001110001111111100000000000000011111111111100000000000000000001000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1031) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000111111111000000000000000000110000001110000000000000000110000000011100000000000000010000000000111000000000000011000000000001000000000000001100000000000000000000000000100001100000000000000000000110011110000000000000000000011111110000000000000000000001111110000000000000000000000111100000000000000000000000111000000000000000000000000011000000000000000000000000011000000000000000000000000011000000000000000000000000011000011110000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1032) begin
            pixels = 784'b0000000000000000000000000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000111100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000001110000000001000000000000000110000001111100000000000000111011111111110000000000000011111111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1033) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000111111110000000000000000011111111111000000000000000111100000100000000000000000110000000000000000000000000011000011000000000000000000011000111100000000000000000001110111100000000000000000000011111000000000000000000000001110000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000001100000011100000000000000001110111111110000000000000000111110001111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1034) begin
            pixels = 784'b0000000000000000000000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000001110000000011100000000000001110000000011110000000000001110000000011110000000000000111110000011110000000000000001111111111110000000000000000000111111110000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1035) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001111110000000000000000000001111111110000000000000000001111111111110000000000000000111100011110000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000001111100000000000000000000000111111000000000000000000000001111100000000000000000000001111100000000000000000000000111100000000000000000000000111100000111000000000000000011110001111100000000000000001110001111100000000000000000111111111100000000000000000011111111100000000000000000000111111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end else if (j == 1036) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111110000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000001000000000000000001111111111111000000000000001111111111111100000000000000111111111000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 1;
        end else if (j == 1037) begin
            pixels = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001111111111000000000000000001111111111110000000000000001111110001111100000000000001111100000011110000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000001111000000000000000000000000111111000000000000000000000001111110000000000000000000000011111000000000000000000000000111100000000000000000000000011100000110000000000000000011111111111000000000000000000111111111100000000000000000011111111110000000000000000000111111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            expected_neuron_out = 2;
        end
    

					 
			#50;
			start = 1;
			#50;
			start = 0;
			
			for (i = 0; i < 810000; i = i + 1) begin
				#50 clk = !clk;
			end clk = 0;

			// update guess count
			if (expected_neuron_out == neuron_out) begin
				guessed_neuron_out = guessed_neuron_out + 1;
			end
		end
	end
endmodule
