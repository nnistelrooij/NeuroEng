module network
#(
	parameter WIDTH = 8,
	parameter HEIGHT = 7,
	// parameter HEIGHT = 784,
	parameter bit [WIDTH:0] WEIGHTS [HEIGHT - 1:0] = '{9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0}
	// parameter bit [WIDTH:0] WEIGHTS [HEIGHT - 1:0] = '{9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0}
)
(
	input wire clk,
	input wire rst,
	input wire [HEIGHT - 1:0] pixels,
	output neuron_out
);
	wire stim;
	reg [HEIGHT - 1:0] pixels_out_pos = 0;
	reg [HEIGHT - 1:0] pixels_out_neg = 0;
	wire [HEIGHT - 1:0] pixels_out;
	wire [HEIGHT - 1:0] tmp;
	
	stim S (
		.clk(clk),
		.rst(rst),
		.stim_out(stim)
	);
	
	genvar i;
	generate
		for (i = 0; i < HEIGHT; i = i + 1) begin : generate_block
			if (WEIGHTS[i][WIDTH]) begin
				divider #(.WIDTH(WIDTH)) Dneg (
					.clk(stim & pixels[i]),
					.rst(rst),
					.w(WEIGHTS[i][WIDTH - 1:0]),
					.neuron_out(pixels_out_neg[i])
				);
			end else begin			
				divider #(.WIDTH(WIDTH)) Dpos (
					.clk(stim & pixels[i]),
					.rst(rst),
					.w(WEIGHTS[i][WIDTH - 1:0]),
					.neuron_out(tmp[i])
				);
				delay De (
					.clk(clk),
					.rst(rst),
					.signal(tmp[i]),
					.neuron_out(pixels_out_pos[i])
				);
			end
		end
	endgenerate

	output2 #(.WIDTH(WIDTH), .HEIGHT(HEIGHT)) Out (
		.clk(clk),
		.rst(rst),
		.inputs(pixels_out),
		.neuron_out(neuron_out)
	);
	
	assign pixels_out = (stim * ~pixels_out_neg) | pixels_out_pos;
endmodule


module testbench_network;
	reg clk = 0;
	reg rst = 1;
	reg [783:0] pixels = 1;
	wire neuron_out;
	
	network #(.HEIGHT(784), .WEIGHTS('{9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0, 9'b0})) N (
		.clk(clk),
		.rst(rst),
		.pixels(pixels),
		.neuron_out(neuron_out)
	);
	
	initial begin
		integer i;
		for (i = 0; i < 1024; i = i + 1) begin
			#50 clk = !clk;
		end
	end
endmodule
